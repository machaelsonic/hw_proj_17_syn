// NIOS2.v

// Generated using ACDS version 12.1 177 at 2017.08.04.17:24:01

`timescale 1 ps / 1 ps
module NIOS2 (
		output wire        epcs_flash_controller_0_external_dclk,    //  epcs_flash_controller_0_external.dclk
		output wire        epcs_flash_controller_0_external_sce,     //                                  .sce
		output wire        epcs_flash_controller_0_external_sdo,     //                                  .sdo
		input  wire        epcs_flash_controller_0_external_data0,   //                                  .data0
		output wire [31:0] tx_data_l_external_connection_export,     //     tx_data_l_external_connection.export
		input  wire        uart_external_connection_rxd,             //          uart_external_connection.rxd
		output wire        uart_external_connection_txd,             //                                  .txd
		output wire        tx_data_valid_external_connection_export, // tx_data_valid_external_connection.export
		input  wire        reset_reset_n,                            //                             reset.reset_n
		input  wire        clk_clk,                                  //                               clk.clk
		input  wire [3:0]  data_external_connection_export,          //          data_external_connection.export
		input  wire        pre_come_external_connection_export,      //      pre_come_external_connection.export
		input  wire [31:0] data_l_external_connection_export,        //        data_l_external_connection.export
		output wire [3:0]  tx_data_h_external_connection_export      //     tx_data_h_external_connection.export
	);

	wire         cpu_instruction_master_waitrequest;                                                                             // CPU_instruction_master_translator:av_waitrequest -> CPU:i_waitrequest
	wire  [18:0] cpu_instruction_master_address;                                                                                 // CPU:i_address -> CPU_instruction_master_translator:av_address
	wire         cpu_instruction_master_read;                                                                                    // CPU:i_read -> CPU_instruction_master_translator:av_read
	wire  [31:0] cpu_instruction_master_readdata;                                                                                // CPU_instruction_master_translator:av_readdata -> CPU:i_readdata
	wire         cpu_instruction_master_readdatavalid;                                                                           // CPU_instruction_master_translator:av_readdatavalid -> CPU:i_readdatavalid
	wire         cpu_data_master_waitrequest;                                                                                    // CPU_data_master_translator:av_waitrequest -> CPU:d_waitrequest
	wire  [31:0] cpu_data_master_writedata;                                                                                      // CPU:d_writedata -> CPU_data_master_translator:av_writedata
	wire  [18:0] cpu_data_master_address;                                                                                        // CPU:d_address -> CPU_data_master_translator:av_address
	wire         cpu_data_master_write;                                                                                          // CPU:d_write -> CPU_data_master_translator:av_write
	wire         cpu_data_master_read;                                                                                           // CPU:d_read -> CPU_data_master_translator:av_read
	wire  [31:0] cpu_data_master_readdata;                                                                                       // CPU_data_master_translator:av_readdata -> CPU:d_readdata
	wire         cpu_data_master_debugaccess;                                                                                    // CPU:jtag_debug_module_debugaccess_to_roms -> CPU_data_master_translator:av_debugaccess
	wire         cpu_data_master_readdatavalid;                                                                                  // CPU_data_master_translator:av_readdatavalid -> CPU:d_readdatavalid
	wire   [3:0] cpu_data_master_byteenable;                                                                                     // CPU:d_byteenable -> CPU_data_master_translator:av_byteenable
	wire  [31:0] cpu_jtag_debug_module_translator_avalon_anti_slave_0_writedata;                                                 // CPU_jtag_debug_module_translator:av_writedata -> CPU:jtag_debug_module_writedata
	wire   [8:0] cpu_jtag_debug_module_translator_avalon_anti_slave_0_address;                                                   // CPU_jtag_debug_module_translator:av_address -> CPU:jtag_debug_module_address
	wire         cpu_jtag_debug_module_translator_avalon_anti_slave_0_chipselect;                                                // CPU_jtag_debug_module_translator:av_chipselect -> CPU:jtag_debug_module_select
	wire         cpu_jtag_debug_module_translator_avalon_anti_slave_0_write;                                                     // CPU_jtag_debug_module_translator:av_write -> CPU:jtag_debug_module_write
	wire  [31:0] cpu_jtag_debug_module_translator_avalon_anti_slave_0_readdata;                                                  // CPU:jtag_debug_module_readdata -> CPU_jtag_debug_module_translator:av_readdata
	wire         cpu_jtag_debug_module_translator_avalon_anti_slave_0_begintransfer;                                             // CPU_jtag_debug_module_translator:av_begintransfer -> CPU:jtag_debug_module_begintransfer
	wire         cpu_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess;                                               // CPU_jtag_debug_module_translator:av_debugaccess -> CPU:jtag_debug_module_debugaccess
	wire   [3:0] cpu_jtag_debug_module_translator_avalon_anti_slave_0_byteenable;                                                // CPU_jtag_debug_module_translator:av_byteenable -> CPU:jtag_debug_module_byteenable
	wire  [31:0] ram_s1_translator_avalon_anti_slave_0_writedata;                                                                // RAM_s1_translator:av_writedata -> RAM:writedata
	wire  [14:0] ram_s1_translator_avalon_anti_slave_0_address;                                                                  // RAM_s1_translator:av_address -> RAM:address
	wire         ram_s1_translator_avalon_anti_slave_0_chipselect;                                                               // RAM_s1_translator:av_chipselect -> RAM:chipselect
	wire         ram_s1_translator_avalon_anti_slave_0_clken;                                                                    // RAM_s1_translator:av_clken -> RAM:clken
	wire         ram_s1_translator_avalon_anti_slave_0_write;                                                                    // RAM_s1_translator:av_write -> RAM:write
	wire  [31:0] ram_s1_translator_avalon_anti_slave_0_readdata;                                                                 // RAM:readdata -> RAM_s1_translator:av_readdata
	wire   [3:0] ram_s1_translator_avalon_anti_slave_0_byteenable;                                                               // RAM_s1_translator:av_byteenable -> RAM:byteenable
	wire  [31:0] epcs_flash_controller_0_epcs_control_port_translator_avalon_anti_slave_0_writedata;                             // epcs_flash_controller_0_epcs_control_port_translator:av_writedata -> epcs_flash_controller_0:writedata
	wire   [8:0] epcs_flash_controller_0_epcs_control_port_translator_avalon_anti_slave_0_address;                               // epcs_flash_controller_0_epcs_control_port_translator:av_address -> epcs_flash_controller_0:address
	wire         epcs_flash_controller_0_epcs_control_port_translator_avalon_anti_slave_0_chipselect;                            // epcs_flash_controller_0_epcs_control_port_translator:av_chipselect -> epcs_flash_controller_0:chipselect
	wire         epcs_flash_controller_0_epcs_control_port_translator_avalon_anti_slave_0_write;                                 // epcs_flash_controller_0_epcs_control_port_translator:av_write -> epcs_flash_controller_0:write_n
	wire         epcs_flash_controller_0_epcs_control_port_translator_avalon_anti_slave_0_read;                                  // epcs_flash_controller_0_epcs_control_port_translator:av_read -> epcs_flash_controller_0:read_n
	wire  [31:0] epcs_flash_controller_0_epcs_control_port_translator_avalon_anti_slave_0_readdata;                              // epcs_flash_controller_0:readdata -> epcs_flash_controller_0_epcs_control_port_translator:av_readdata
	wire  [15:0] uart_s1_translator_avalon_anti_slave_0_writedata;                                                               // uart_s1_translator:av_writedata -> uart:writedata
	wire   [2:0] uart_s1_translator_avalon_anti_slave_0_address;                                                                 // uart_s1_translator:av_address -> uart:address
	wire         uart_s1_translator_avalon_anti_slave_0_chipselect;                                                              // uart_s1_translator:av_chipselect -> uart:chipselect
	wire         uart_s1_translator_avalon_anti_slave_0_write;                                                                   // uart_s1_translator:av_write -> uart:write_n
	wire         uart_s1_translator_avalon_anti_slave_0_read;                                                                    // uart_s1_translator:av_read -> uart:read_n
	wire  [15:0] uart_s1_translator_avalon_anti_slave_0_readdata;                                                                // uart:readdata -> uart_s1_translator:av_readdata
	wire         uart_s1_translator_avalon_anti_slave_0_begintransfer;                                                           // uart_s1_translator:av_begintransfer -> uart:begintransfer
	wire         jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest;                                         // jtag_uart:av_waitrequest -> jtag_uart_avalon_jtag_slave_translator:av_waitrequest
	wire  [31:0] jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata;                                           // jtag_uart_avalon_jtag_slave_translator:av_writedata -> jtag_uart:av_writedata
	wire   [0:0] jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_address;                                             // jtag_uart_avalon_jtag_slave_translator:av_address -> jtag_uart:av_address
	wire         jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect;                                          // jtag_uart_avalon_jtag_slave_translator:av_chipselect -> jtag_uart:av_chipselect
	wire         jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_write;                                               // jtag_uart_avalon_jtag_slave_translator:av_write -> jtag_uart:av_write_n
	wire         jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_read;                                                // jtag_uart_avalon_jtag_slave_translator:av_read -> jtag_uart:av_read_n
	wire  [31:0] jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata;                                            // jtag_uart:av_readdata -> jtag_uart_avalon_jtag_slave_translator:av_readdata
	wire   [1:0] data_h_s1_translator_avalon_anti_slave_0_address;                                                               // DATA_H_s1_translator:av_address -> DATA_H:address
	wire  [31:0] data_h_s1_translator_avalon_anti_slave_0_readdata;                                                              // DATA_H:readdata -> DATA_H_s1_translator:av_readdata
	wire   [0:0] sysid_control_slave_translator_avalon_anti_slave_0_address;                                                     // sysid_control_slave_translator:av_address -> sysid:address
	wire  [31:0] sysid_control_slave_translator_avalon_anti_slave_0_readdata;                                                    // sysid:readdata -> sysid_control_slave_translator:av_readdata
	wire   [1:0] data_l_s1_translator_avalon_anti_slave_0_address;                                                               // DATA_L_s1_translator:av_address -> DATA_L:address
	wire  [31:0] data_l_s1_translator_avalon_anti_slave_0_readdata;                                                              // DATA_L:readdata -> DATA_L_s1_translator:av_readdata
	wire  [31:0] pre_come_s1_translator_avalon_anti_slave_0_writedata;                                                           // pre_come_s1_translator:av_writedata -> pre_come:writedata
	wire   [1:0] pre_come_s1_translator_avalon_anti_slave_0_address;                                                             // pre_come_s1_translator:av_address -> pre_come:address
	wire         pre_come_s1_translator_avalon_anti_slave_0_chipselect;                                                          // pre_come_s1_translator:av_chipselect -> pre_come:chipselect
	wire         pre_come_s1_translator_avalon_anti_slave_0_write;                                                               // pre_come_s1_translator:av_write -> pre_come:write_n
	wire  [31:0] pre_come_s1_translator_avalon_anti_slave_0_readdata;                                                            // pre_come:readdata -> pre_come_s1_translator:av_readdata
	wire  [31:0] tx_data_l_s1_translator_avalon_anti_slave_0_writedata;                                                          // TX_DATA_L_s1_translator:av_writedata -> TX_DATA_L:writedata
	wire   [1:0] tx_data_l_s1_translator_avalon_anti_slave_0_address;                                                            // TX_DATA_L_s1_translator:av_address -> TX_DATA_L:address
	wire         tx_data_l_s1_translator_avalon_anti_slave_0_chipselect;                                                         // TX_DATA_L_s1_translator:av_chipselect -> TX_DATA_L:chipselect
	wire         tx_data_l_s1_translator_avalon_anti_slave_0_write;                                                              // TX_DATA_L_s1_translator:av_write -> TX_DATA_L:write_n
	wire  [31:0] tx_data_l_s1_translator_avalon_anti_slave_0_readdata;                                                           // TX_DATA_L:readdata -> TX_DATA_L_s1_translator:av_readdata
	wire  [31:0] tx_data_h_s1_translator_avalon_anti_slave_0_writedata;                                                          // TX_DATA_H_s1_translator:av_writedata -> TX_DATA_H:writedata
	wire   [1:0] tx_data_h_s1_translator_avalon_anti_slave_0_address;                                                            // TX_DATA_H_s1_translator:av_address -> TX_DATA_H:address
	wire         tx_data_h_s1_translator_avalon_anti_slave_0_chipselect;                                                         // TX_DATA_H_s1_translator:av_chipselect -> TX_DATA_H:chipselect
	wire         tx_data_h_s1_translator_avalon_anti_slave_0_write;                                                              // TX_DATA_H_s1_translator:av_write -> TX_DATA_H:write_n
	wire  [31:0] tx_data_h_s1_translator_avalon_anti_slave_0_readdata;                                                           // TX_DATA_H:readdata -> TX_DATA_H_s1_translator:av_readdata
	wire  [31:0] tx_data_valid_s1_translator_avalon_anti_slave_0_writedata;                                                      // TX_DATA_VALID_s1_translator:av_writedata -> TX_DATA_VALID:writedata
	wire   [1:0] tx_data_valid_s1_translator_avalon_anti_slave_0_address;                                                        // TX_DATA_VALID_s1_translator:av_address -> TX_DATA_VALID:address
	wire         tx_data_valid_s1_translator_avalon_anti_slave_0_chipselect;                                                     // TX_DATA_VALID_s1_translator:av_chipselect -> TX_DATA_VALID:chipselect
	wire         tx_data_valid_s1_translator_avalon_anti_slave_0_write;                                                          // TX_DATA_VALID_s1_translator:av_write -> TX_DATA_VALID:write_n
	wire  [31:0] tx_data_valid_s1_translator_avalon_anti_slave_0_readdata;                                                       // TX_DATA_VALID:readdata -> TX_DATA_VALID_s1_translator:av_readdata
	wire         cpu_instruction_master_translator_avalon_universal_master_0_waitrequest;                                        // CPU_instruction_master_translator_avalon_universal_master_0_agent:av_waitrequest -> CPU_instruction_master_translator:uav_waitrequest
	wire   [2:0] cpu_instruction_master_translator_avalon_universal_master_0_burstcount;                                         // CPU_instruction_master_translator:uav_burstcount -> CPU_instruction_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire  [31:0] cpu_instruction_master_translator_avalon_universal_master_0_writedata;                                          // CPU_instruction_master_translator:uav_writedata -> CPU_instruction_master_translator_avalon_universal_master_0_agent:av_writedata
	wire  [18:0] cpu_instruction_master_translator_avalon_universal_master_0_address;                                            // CPU_instruction_master_translator:uav_address -> CPU_instruction_master_translator_avalon_universal_master_0_agent:av_address
	wire         cpu_instruction_master_translator_avalon_universal_master_0_lock;                                               // CPU_instruction_master_translator:uav_lock -> CPU_instruction_master_translator_avalon_universal_master_0_agent:av_lock
	wire         cpu_instruction_master_translator_avalon_universal_master_0_write;                                              // CPU_instruction_master_translator:uav_write -> CPU_instruction_master_translator_avalon_universal_master_0_agent:av_write
	wire         cpu_instruction_master_translator_avalon_universal_master_0_read;                                               // CPU_instruction_master_translator:uav_read -> CPU_instruction_master_translator_avalon_universal_master_0_agent:av_read
	wire  [31:0] cpu_instruction_master_translator_avalon_universal_master_0_readdata;                                           // CPU_instruction_master_translator_avalon_universal_master_0_agent:av_readdata -> CPU_instruction_master_translator:uav_readdata
	wire         cpu_instruction_master_translator_avalon_universal_master_0_debugaccess;                                        // CPU_instruction_master_translator:uav_debugaccess -> CPU_instruction_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire   [3:0] cpu_instruction_master_translator_avalon_universal_master_0_byteenable;                                         // CPU_instruction_master_translator:uav_byteenable -> CPU_instruction_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire         cpu_instruction_master_translator_avalon_universal_master_0_readdatavalid;                                      // CPU_instruction_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> CPU_instruction_master_translator:uav_readdatavalid
	wire         cpu_data_master_translator_avalon_universal_master_0_waitrequest;                                               // CPU_data_master_translator_avalon_universal_master_0_agent:av_waitrequest -> CPU_data_master_translator:uav_waitrequest
	wire   [2:0] cpu_data_master_translator_avalon_universal_master_0_burstcount;                                                // CPU_data_master_translator:uav_burstcount -> CPU_data_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire  [31:0] cpu_data_master_translator_avalon_universal_master_0_writedata;                                                 // CPU_data_master_translator:uav_writedata -> CPU_data_master_translator_avalon_universal_master_0_agent:av_writedata
	wire  [18:0] cpu_data_master_translator_avalon_universal_master_0_address;                                                   // CPU_data_master_translator:uav_address -> CPU_data_master_translator_avalon_universal_master_0_agent:av_address
	wire         cpu_data_master_translator_avalon_universal_master_0_lock;                                                      // CPU_data_master_translator:uav_lock -> CPU_data_master_translator_avalon_universal_master_0_agent:av_lock
	wire         cpu_data_master_translator_avalon_universal_master_0_write;                                                     // CPU_data_master_translator:uav_write -> CPU_data_master_translator_avalon_universal_master_0_agent:av_write
	wire         cpu_data_master_translator_avalon_universal_master_0_read;                                                      // CPU_data_master_translator:uav_read -> CPU_data_master_translator_avalon_universal_master_0_agent:av_read
	wire  [31:0] cpu_data_master_translator_avalon_universal_master_0_readdata;                                                  // CPU_data_master_translator_avalon_universal_master_0_agent:av_readdata -> CPU_data_master_translator:uav_readdata
	wire         cpu_data_master_translator_avalon_universal_master_0_debugaccess;                                               // CPU_data_master_translator:uav_debugaccess -> CPU_data_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire   [3:0] cpu_data_master_translator_avalon_universal_master_0_byteenable;                                                // CPU_data_master_translator:uav_byteenable -> CPU_data_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire         cpu_data_master_translator_avalon_universal_master_0_readdatavalid;                                             // CPU_data_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> CPU_data_master_translator:uav_readdatavalid
	wire         cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                 // CPU_jtag_debug_module_translator:uav_waitrequest -> CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount;                                  // CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_burstcount -> CPU_jtag_debug_module_translator:uav_burstcount
	wire  [31:0] cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata;                                   // CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_writedata -> CPU_jtag_debug_module_translator:uav_writedata
	wire  [18:0] cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address;                                     // CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_address -> CPU_jtag_debug_module_translator:uav_address
	wire         cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write;                                       // CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_write -> CPU_jtag_debug_module_translator:uav_write
	wire         cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock;                                        // CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_lock -> CPU_jtag_debug_module_translator:uav_lock
	wire         cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read;                                        // CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_read -> CPU_jtag_debug_module_translator:uav_read
	wire  [31:0] cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata;                                    // CPU_jtag_debug_module_translator:uav_readdata -> CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                               // CPU_jtag_debug_module_translator:uav_readdatavalid -> CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                 // CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_debugaccess -> CPU_jtag_debug_module_translator:uav_debugaccess
	wire   [3:0] cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable;                                  // CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_byteenable -> CPU_jtag_debug_module_translator:uav_byteenable
	wire         cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                          // CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid;                                // CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_valid -> CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                        // CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [94:0] cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data;                                 // CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_data -> CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready;                                // CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                       // CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                             // CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                     // CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [94:0] cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                              // CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                             // CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_ready -> CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                           // CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                            // CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                           // CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         ram_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                                // RAM_s1_translator:uav_waitrequest -> RAM_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] ram_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                                 // RAM_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> RAM_s1_translator:uav_burstcount
	wire  [31:0] ram_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                                  // RAM_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> RAM_s1_translator:uav_writedata
	wire  [18:0] ram_s1_translator_avalon_universal_slave_0_agent_m0_address;                                                    // RAM_s1_translator_avalon_universal_slave_0_agent:m0_address -> RAM_s1_translator:uav_address
	wire         ram_s1_translator_avalon_universal_slave_0_agent_m0_write;                                                      // RAM_s1_translator_avalon_universal_slave_0_agent:m0_write -> RAM_s1_translator:uav_write
	wire         ram_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                                       // RAM_s1_translator_avalon_universal_slave_0_agent:m0_lock -> RAM_s1_translator:uav_lock
	wire         ram_s1_translator_avalon_universal_slave_0_agent_m0_read;                                                       // RAM_s1_translator_avalon_universal_slave_0_agent:m0_read -> RAM_s1_translator:uav_read
	wire  [31:0] ram_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                                   // RAM_s1_translator:uav_readdata -> RAM_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         ram_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                              // RAM_s1_translator:uav_readdatavalid -> RAM_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         ram_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                                // RAM_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> RAM_s1_translator:uav_debugaccess
	wire   [3:0] ram_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                                 // RAM_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> RAM_s1_translator:uav_byteenable
	wire         ram_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                                         // RAM_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> RAM_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         ram_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                               // RAM_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> RAM_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         ram_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                                       // RAM_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> RAM_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [94:0] ram_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                                // RAM_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> RAM_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         ram_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                               // RAM_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> RAM_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                                      // RAM_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> RAM_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                            // RAM_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> RAM_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                                    // RAM_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> RAM_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [94:0] ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                             // RAM_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> RAM_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                            // RAM_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> RAM_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         ram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                                          // RAM_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> RAM_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] ram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                           // RAM_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> RAM_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         ram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                                          // RAM_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> RAM_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_waitrequest;             // epcs_flash_controller_0_epcs_control_port_translator:uav_waitrequest -> epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_burstcount;              // epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent:m0_burstcount -> epcs_flash_controller_0_epcs_control_port_translator:uav_burstcount
	wire  [31:0] epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_writedata;               // epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent:m0_writedata -> epcs_flash_controller_0_epcs_control_port_translator:uav_writedata
	wire  [18:0] epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_address;                 // epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent:m0_address -> epcs_flash_controller_0_epcs_control_port_translator:uav_address
	wire         epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_write;                   // epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent:m0_write -> epcs_flash_controller_0_epcs_control_port_translator:uav_write
	wire         epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_lock;                    // epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent:m0_lock -> epcs_flash_controller_0_epcs_control_port_translator:uav_lock
	wire         epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_read;                    // epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent:m0_read -> epcs_flash_controller_0_epcs_control_port_translator:uav_read
	wire  [31:0] epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_readdata;                // epcs_flash_controller_0_epcs_control_port_translator:uav_readdata -> epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_readdatavalid;           // epcs_flash_controller_0_epcs_control_port_translator:uav_readdatavalid -> epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_debugaccess;             // epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent:m0_debugaccess -> epcs_flash_controller_0_epcs_control_port_translator:uav_debugaccess
	wire   [3:0] epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_byteenable;              // epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent:m0_byteenable -> epcs_flash_controller_0_epcs_control_port_translator:uav_byteenable
	wire         epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;      // epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_rf_source_valid;            // epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent:rf_source_valid -> epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;    // epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [94:0] epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_rf_source_data;             // epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent:rf_source_data -> epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_rf_source_ready;            // epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;   // epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;         // epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket; // epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [94:0] epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;          // epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;         // epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent:rf_sink_ready -> epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;       // epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;        // epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;       // epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         uart_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                               // uart_s1_translator:uav_waitrequest -> uart_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] uart_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                                // uart_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> uart_s1_translator:uav_burstcount
	wire  [31:0] uart_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                                 // uart_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> uart_s1_translator:uav_writedata
	wire  [18:0] uart_s1_translator_avalon_universal_slave_0_agent_m0_address;                                                   // uart_s1_translator_avalon_universal_slave_0_agent:m0_address -> uart_s1_translator:uav_address
	wire         uart_s1_translator_avalon_universal_slave_0_agent_m0_write;                                                     // uart_s1_translator_avalon_universal_slave_0_agent:m0_write -> uart_s1_translator:uav_write
	wire         uart_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                                      // uart_s1_translator_avalon_universal_slave_0_agent:m0_lock -> uart_s1_translator:uav_lock
	wire         uart_s1_translator_avalon_universal_slave_0_agent_m0_read;                                                      // uart_s1_translator_avalon_universal_slave_0_agent:m0_read -> uart_s1_translator:uav_read
	wire  [31:0] uart_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                                  // uart_s1_translator:uav_readdata -> uart_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         uart_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                             // uart_s1_translator:uav_readdatavalid -> uart_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         uart_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                               // uart_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> uart_s1_translator:uav_debugaccess
	wire   [3:0] uart_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                                // uart_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> uart_s1_translator:uav_byteenable
	wire         uart_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                                        // uart_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> uart_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         uart_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                              // uart_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> uart_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         uart_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                                      // uart_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> uart_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [94:0] uart_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                               // uart_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> uart_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         uart_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                              // uart_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> uart_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         uart_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                                     // uart_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> uart_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         uart_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                           // uart_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> uart_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         uart_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                                   // uart_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> uart_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [94:0] uart_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                            // uart_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> uart_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         uart_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                           // uart_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> uart_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         uart_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                                         // uart_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> uart_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] uart_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                          // uart_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> uart_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         uart_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                                         // uart_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> uart_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;                           // jtag_uart_avalon_jtag_slave_translator:uav_waitrequest -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                            // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> jtag_uart_avalon_jtag_slave_translator:uav_burstcount
	wire  [31:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                             // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> jtag_uart_avalon_jtag_slave_translator:uav_writedata
	wire  [18:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address;                               // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_address -> jtag_uart_avalon_jtag_slave_translator:uav_address
	wire         jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write;                                 // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_write -> jtag_uart_avalon_jtag_slave_translator:uav_write
	wire         jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock;                                  // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_lock -> jtag_uart_avalon_jtag_slave_translator:uav_lock
	wire         jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read;                                  // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_read -> jtag_uart_avalon_jtag_slave_translator:uav_read
	wire  [31:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                              // jtag_uart_avalon_jtag_slave_translator:uav_readdata -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                         // jtag_uart_avalon_jtag_slave_translator:uav_readdatavalid -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;                           // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> jtag_uart_avalon_jtag_slave_translator:uav_debugaccess
	wire   [3:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                            // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> jtag_uart_avalon_jtag_slave_translator:uav_byteenable
	wire         jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                    // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;                          // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                  // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [94:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data;                           // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;                          // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                 // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                       // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;               // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [94:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                        // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                       // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                     // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                      // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                     // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         data_h_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                             // DATA_H_s1_translator:uav_waitrequest -> DATA_H_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] data_h_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                              // DATA_H_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> DATA_H_s1_translator:uav_burstcount
	wire  [31:0] data_h_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                               // DATA_H_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> DATA_H_s1_translator:uav_writedata
	wire  [18:0] data_h_s1_translator_avalon_universal_slave_0_agent_m0_address;                                                 // DATA_H_s1_translator_avalon_universal_slave_0_agent:m0_address -> DATA_H_s1_translator:uav_address
	wire         data_h_s1_translator_avalon_universal_slave_0_agent_m0_write;                                                   // DATA_H_s1_translator_avalon_universal_slave_0_agent:m0_write -> DATA_H_s1_translator:uav_write
	wire         data_h_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                                    // DATA_H_s1_translator_avalon_universal_slave_0_agent:m0_lock -> DATA_H_s1_translator:uav_lock
	wire         data_h_s1_translator_avalon_universal_slave_0_agent_m0_read;                                                    // DATA_H_s1_translator_avalon_universal_slave_0_agent:m0_read -> DATA_H_s1_translator:uav_read
	wire  [31:0] data_h_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                                // DATA_H_s1_translator:uav_readdata -> DATA_H_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         data_h_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                           // DATA_H_s1_translator:uav_readdatavalid -> DATA_H_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         data_h_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                             // DATA_H_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> DATA_H_s1_translator:uav_debugaccess
	wire   [3:0] data_h_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                              // DATA_H_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> DATA_H_s1_translator:uav_byteenable
	wire         data_h_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                                      // DATA_H_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> DATA_H_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         data_h_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                            // DATA_H_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> DATA_H_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         data_h_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                                    // DATA_H_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> DATA_H_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [94:0] data_h_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                             // DATA_H_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> DATA_H_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         data_h_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                            // DATA_H_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> DATA_H_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         data_h_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                                   // DATA_H_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> DATA_H_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         data_h_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                         // DATA_H_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> DATA_H_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         data_h_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                                 // DATA_H_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> DATA_H_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [94:0] data_h_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                          // DATA_H_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> DATA_H_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         data_h_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                         // DATA_H_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> DATA_H_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         data_h_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                                       // DATA_H_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> DATA_H_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] data_h_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                        // DATA_H_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> DATA_H_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         data_h_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                                       // DATA_H_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> DATA_H_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                   // sysid_control_slave_translator:uav_waitrequest -> sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                                    // sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> sysid_control_slave_translator:uav_burstcount
	wire  [31:0] sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                                     // sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> sysid_control_slave_translator:uav_writedata
	wire  [18:0] sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_address;                                       // sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_address -> sysid_control_slave_translator:uav_address
	wire         sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_write;                                         // sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_write -> sysid_control_slave_translator:uav_write
	wire         sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_lock;                                          // sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_lock -> sysid_control_slave_translator:uav_lock
	wire         sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_read;                                          // sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_read -> sysid_control_slave_translator:uav_read
	wire  [31:0] sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                                      // sysid_control_slave_translator:uav_readdata -> sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                 // sysid_control_slave_translator:uav_readdatavalid -> sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                   // sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> sysid_control_slave_translator:uav_debugaccess
	wire   [3:0] sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                                    // sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> sysid_control_slave_translator:uav_byteenable
	wire         sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                            // sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;                                  // sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                          // sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [94:0] sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data;                                   // sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;                                  // sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                         // sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                               // sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                       // sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [94:0] sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                // sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                               // sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                             // sysid_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                              // sysid_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                             // sysid_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         data_l_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                             // DATA_L_s1_translator:uav_waitrequest -> DATA_L_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] data_l_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                              // DATA_L_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> DATA_L_s1_translator:uav_burstcount
	wire  [31:0] data_l_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                               // DATA_L_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> DATA_L_s1_translator:uav_writedata
	wire  [18:0] data_l_s1_translator_avalon_universal_slave_0_agent_m0_address;                                                 // DATA_L_s1_translator_avalon_universal_slave_0_agent:m0_address -> DATA_L_s1_translator:uav_address
	wire         data_l_s1_translator_avalon_universal_slave_0_agent_m0_write;                                                   // DATA_L_s1_translator_avalon_universal_slave_0_agent:m0_write -> DATA_L_s1_translator:uav_write
	wire         data_l_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                                    // DATA_L_s1_translator_avalon_universal_slave_0_agent:m0_lock -> DATA_L_s1_translator:uav_lock
	wire         data_l_s1_translator_avalon_universal_slave_0_agent_m0_read;                                                    // DATA_L_s1_translator_avalon_universal_slave_0_agent:m0_read -> DATA_L_s1_translator:uav_read
	wire  [31:0] data_l_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                                // DATA_L_s1_translator:uav_readdata -> DATA_L_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         data_l_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                           // DATA_L_s1_translator:uav_readdatavalid -> DATA_L_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         data_l_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                             // DATA_L_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> DATA_L_s1_translator:uav_debugaccess
	wire   [3:0] data_l_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                              // DATA_L_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> DATA_L_s1_translator:uav_byteenable
	wire         data_l_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                                      // DATA_L_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> DATA_L_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         data_l_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                            // DATA_L_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> DATA_L_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         data_l_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                                    // DATA_L_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> DATA_L_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [94:0] data_l_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                             // DATA_L_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> DATA_L_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         data_l_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                            // DATA_L_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> DATA_L_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         data_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                                   // DATA_L_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> DATA_L_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         data_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                         // DATA_L_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> DATA_L_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         data_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                                 // DATA_L_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> DATA_L_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [94:0] data_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                          // DATA_L_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> DATA_L_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         data_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                         // DATA_L_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> DATA_L_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         data_l_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                                       // DATA_L_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> DATA_L_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] data_l_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                        // DATA_L_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> DATA_L_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         data_l_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                                       // DATA_L_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> DATA_L_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         pre_come_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                           // pre_come_s1_translator:uav_waitrequest -> pre_come_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] pre_come_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                            // pre_come_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> pre_come_s1_translator:uav_burstcount
	wire  [31:0] pre_come_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                             // pre_come_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> pre_come_s1_translator:uav_writedata
	wire  [18:0] pre_come_s1_translator_avalon_universal_slave_0_agent_m0_address;                                               // pre_come_s1_translator_avalon_universal_slave_0_agent:m0_address -> pre_come_s1_translator:uav_address
	wire         pre_come_s1_translator_avalon_universal_slave_0_agent_m0_write;                                                 // pre_come_s1_translator_avalon_universal_slave_0_agent:m0_write -> pre_come_s1_translator:uav_write
	wire         pre_come_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                                  // pre_come_s1_translator_avalon_universal_slave_0_agent:m0_lock -> pre_come_s1_translator:uav_lock
	wire         pre_come_s1_translator_avalon_universal_slave_0_agent_m0_read;                                                  // pre_come_s1_translator_avalon_universal_slave_0_agent:m0_read -> pre_come_s1_translator:uav_read
	wire  [31:0] pre_come_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                              // pre_come_s1_translator:uav_readdata -> pre_come_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         pre_come_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                         // pre_come_s1_translator:uav_readdatavalid -> pre_come_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         pre_come_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                           // pre_come_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> pre_come_s1_translator:uav_debugaccess
	wire   [3:0] pre_come_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                            // pre_come_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> pre_come_s1_translator:uav_byteenable
	wire         pre_come_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                                    // pre_come_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> pre_come_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         pre_come_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                          // pre_come_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> pre_come_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         pre_come_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                                  // pre_come_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> pre_come_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [94:0] pre_come_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                           // pre_come_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> pre_come_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         pre_come_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                          // pre_come_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> pre_come_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         pre_come_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                                 // pre_come_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> pre_come_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         pre_come_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                       // pre_come_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> pre_come_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         pre_come_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                               // pre_come_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> pre_come_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [94:0] pre_come_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                        // pre_come_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> pre_come_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         pre_come_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                       // pre_come_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> pre_come_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         pre_come_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                                     // pre_come_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> pre_come_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] pre_come_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                      // pre_come_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> pre_come_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         pre_come_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                                     // pre_come_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> pre_come_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         tx_data_l_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                          // TX_DATA_L_s1_translator:uav_waitrequest -> TX_DATA_L_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] tx_data_l_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                           // TX_DATA_L_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> TX_DATA_L_s1_translator:uav_burstcount
	wire  [31:0] tx_data_l_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                            // TX_DATA_L_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> TX_DATA_L_s1_translator:uav_writedata
	wire  [18:0] tx_data_l_s1_translator_avalon_universal_slave_0_agent_m0_address;                                              // TX_DATA_L_s1_translator_avalon_universal_slave_0_agent:m0_address -> TX_DATA_L_s1_translator:uav_address
	wire         tx_data_l_s1_translator_avalon_universal_slave_0_agent_m0_write;                                                // TX_DATA_L_s1_translator_avalon_universal_slave_0_agent:m0_write -> TX_DATA_L_s1_translator:uav_write
	wire         tx_data_l_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                                 // TX_DATA_L_s1_translator_avalon_universal_slave_0_agent:m0_lock -> TX_DATA_L_s1_translator:uav_lock
	wire         tx_data_l_s1_translator_avalon_universal_slave_0_agent_m0_read;                                                 // TX_DATA_L_s1_translator_avalon_universal_slave_0_agent:m0_read -> TX_DATA_L_s1_translator:uav_read
	wire  [31:0] tx_data_l_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                             // TX_DATA_L_s1_translator:uav_readdata -> TX_DATA_L_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         tx_data_l_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                        // TX_DATA_L_s1_translator:uav_readdatavalid -> TX_DATA_L_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         tx_data_l_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                          // TX_DATA_L_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> TX_DATA_L_s1_translator:uav_debugaccess
	wire   [3:0] tx_data_l_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                           // TX_DATA_L_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> TX_DATA_L_s1_translator:uav_byteenable
	wire         tx_data_l_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                                   // TX_DATA_L_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> TX_DATA_L_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         tx_data_l_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                         // TX_DATA_L_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> TX_DATA_L_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         tx_data_l_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                                 // TX_DATA_L_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> TX_DATA_L_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [94:0] tx_data_l_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                          // TX_DATA_L_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> TX_DATA_L_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         tx_data_l_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                         // TX_DATA_L_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> TX_DATA_L_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         tx_data_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                                // TX_DATA_L_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> TX_DATA_L_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         tx_data_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                      // TX_DATA_L_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> TX_DATA_L_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         tx_data_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                              // TX_DATA_L_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> TX_DATA_L_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [94:0] tx_data_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                       // TX_DATA_L_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> TX_DATA_L_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         tx_data_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                      // TX_DATA_L_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> TX_DATA_L_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         tx_data_l_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                                    // TX_DATA_L_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> TX_DATA_L_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] tx_data_l_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                     // TX_DATA_L_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> TX_DATA_L_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         tx_data_l_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                                    // TX_DATA_L_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> TX_DATA_L_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         tx_data_h_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                          // TX_DATA_H_s1_translator:uav_waitrequest -> TX_DATA_H_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] tx_data_h_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                           // TX_DATA_H_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> TX_DATA_H_s1_translator:uav_burstcount
	wire  [31:0] tx_data_h_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                            // TX_DATA_H_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> TX_DATA_H_s1_translator:uav_writedata
	wire  [18:0] tx_data_h_s1_translator_avalon_universal_slave_0_agent_m0_address;                                              // TX_DATA_H_s1_translator_avalon_universal_slave_0_agent:m0_address -> TX_DATA_H_s1_translator:uav_address
	wire         tx_data_h_s1_translator_avalon_universal_slave_0_agent_m0_write;                                                // TX_DATA_H_s1_translator_avalon_universal_slave_0_agent:m0_write -> TX_DATA_H_s1_translator:uav_write
	wire         tx_data_h_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                                 // TX_DATA_H_s1_translator_avalon_universal_slave_0_agent:m0_lock -> TX_DATA_H_s1_translator:uav_lock
	wire         tx_data_h_s1_translator_avalon_universal_slave_0_agent_m0_read;                                                 // TX_DATA_H_s1_translator_avalon_universal_slave_0_agent:m0_read -> TX_DATA_H_s1_translator:uav_read
	wire  [31:0] tx_data_h_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                             // TX_DATA_H_s1_translator:uav_readdata -> TX_DATA_H_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         tx_data_h_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                        // TX_DATA_H_s1_translator:uav_readdatavalid -> TX_DATA_H_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         tx_data_h_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                          // TX_DATA_H_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> TX_DATA_H_s1_translator:uav_debugaccess
	wire   [3:0] tx_data_h_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                           // TX_DATA_H_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> TX_DATA_H_s1_translator:uav_byteenable
	wire         tx_data_h_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                                   // TX_DATA_H_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> TX_DATA_H_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         tx_data_h_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                         // TX_DATA_H_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> TX_DATA_H_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         tx_data_h_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                                 // TX_DATA_H_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> TX_DATA_H_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [94:0] tx_data_h_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                          // TX_DATA_H_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> TX_DATA_H_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         tx_data_h_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                         // TX_DATA_H_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> TX_DATA_H_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         tx_data_h_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                                // TX_DATA_H_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> TX_DATA_H_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         tx_data_h_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                      // TX_DATA_H_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> TX_DATA_H_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         tx_data_h_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                              // TX_DATA_H_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> TX_DATA_H_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [94:0] tx_data_h_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                       // TX_DATA_H_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> TX_DATA_H_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         tx_data_h_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                      // TX_DATA_H_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> TX_DATA_H_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         tx_data_h_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                                    // TX_DATA_H_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> TX_DATA_H_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] tx_data_h_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                     // TX_DATA_H_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> TX_DATA_H_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         tx_data_h_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                                    // TX_DATA_H_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> TX_DATA_H_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         tx_data_valid_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                      // TX_DATA_VALID_s1_translator:uav_waitrequest -> TX_DATA_VALID_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] tx_data_valid_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                       // TX_DATA_VALID_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> TX_DATA_VALID_s1_translator:uav_burstcount
	wire  [31:0] tx_data_valid_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                        // TX_DATA_VALID_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> TX_DATA_VALID_s1_translator:uav_writedata
	wire  [18:0] tx_data_valid_s1_translator_avalon_universal_slave_0_agent_m0_address;                                          // TX_DATA_VALID_s1_translator_avalon_universal_slave_0_agent:m0_address -> TX_DATA_VALID_s1_translator:uav_address
	wire         tx_data_valid_s1_translator_avalon_universal_slave_0_agent_m0_write;                                            // TX_DATA_VALID_s1_translator_avalon_universal_slave_0_agent:m0_write -> TX_DATA_VALID_s1_translator:uav_write
	wire         tx_data_valid_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                             // TX_DATA_VALID_s1_translator_avalon_universal_slave_0_agent:m0_lock -> TX_DATA_VALID_s1_translator:uav_lock
	wire         tx_data_valid_s1_translator_avalon_universal_slave_0_agent_m0_read;                                             // TX_DATA_VALID_s1_translator_avalon_universal_slave_0_agent:m0_read -> TX_DATA_VALID_s1_translator:uav_read
	wire  [31:0] tx_data_valid_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                         // TX_DATA_VALID_s1_translator:uav_readdata -> TX_DATA_VALID_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         tx_data_valid_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                    // TX_DATA_VALID_s1_translator:uav_readdatavalid -> TX_DATA_VALID_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         tx_data_valid_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                      // TX_DATA_VALID_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> TX_DATA_VALID_s1_translator:uav_debugaccess
	wire   [3:0] tx_data_valid_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                       // TX_DATA_VALID_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> TX_DATA_VALID_s1_translator:uav_byteenable
	wire         tx_data_valid_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                               // TX_DATA_VALID_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> TX_DATA_VALID_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         tx_data_valid_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                     // TX_DATA_VALID_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> TX_DATA_VALID_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         tx_data_valid_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                             // TX_DATA_VALID_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> TX_DATA_VALID_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [94:0] tx_data_valid_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                      // TX_DATA_VALID_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> TX_DATA_VALID_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         tx_data_valid_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                     // TX_DATA_VALID_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> TX_DATA_VALID_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         tx_data_valid_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                            // TX_DATA_VALID_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> TX_DATA_VALID_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         tx_data_valid_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                  // TX_DATA_VALID_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> TX_DATA_VALID_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         tx_data_valid_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                          // TX_DATA_VALID_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> TX_DATA_VALID_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [94:0] tx_data_valid_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                   // TX_DATA_VALID_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> TX_DATA_VALID_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         tx_data_valid_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                  // TX_DATA_VALID_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> TX_DATA_VALID_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         tx_data_valid_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                                // TX_DATA_VALID_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> TX_DATA_VALID_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] tx_data_valid_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                 // TX_DATA_VALID_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> TX_DATA_VALID_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         tx_data_valid_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                                // TX_DATA_VALID_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> TX_DATA_VALID_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket;                               // CPU_instruction_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router:sink_endofpacket
	wire         cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_valid;                                     // CPU_instruction_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router:sink_valid
	wire         cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket;                             // CPU_instruction_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router:sink_startofpacket
	wire  [93:0] cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_data;                                      // CPU_instruction_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router:sink_data
	wire         cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_ready;                                     // addr_router:sink_ready -> CPU_instruction_master_translator_avalon_universal_master_0_agent:cp_ready
	wire         cpu_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket;                                      // CPU_data_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_001:sink_endofpacket
	wire         cpu_data_master_translator_avalon_universal_master_0_agent_cp_valid;                                            // CPU_data_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_001:sink_valid
	wire         cpu_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket;                                    // CPU_data_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_001:sink_startofpacket
	wire  [93:0] cpu_data_master_translator_avalon_universal_master_0_agent_cp_data;                                             // CPU_data_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router_001:sink_data
	wire         cpu_data_master_translator_avalon_universal_master_0_agent_cp_ready;                                            // addr_router_001:sink_ready -> CPU_data_master_translator_avalon_universal_master_0_agent:cp_ready
	wire         cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                 // CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router:sink_endofpacket
	wire         cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid;                                       // CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_valid -> id_router:sink_valid
	wire         cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket;                               // CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router:sink_startofpacket
	wire  [93:0] cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data;                                        // CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_data -> id_router:sink_data
	wire         cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready;                                       // id_router:sink_ready -> CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_ready
	wire         ram_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                                // RAM_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_001:sink_endofpacket
	wire         ram_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                                      // RAM_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_001:sink_valid
	wire         ram_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                              // RAM_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_001:sink_startofpacket
	wire  [93:0] ram_s1_translator_avalon_universal_slave_0_agent_rp_data;                                                       // RAM_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_001:sink_data
	wire         ram_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                                      // id_router_001:sink_ready -> RAM_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_rp_endofpacket;             // epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_002:sink_endofpacket
	wire         epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_rp_valid;                   // epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_002:sink_valid
	wire         epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_rp_startofpacket;           // epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_002:sink_startofpacket
	wire  [93:0] epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_rp_data;                    // epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent:rp_data -> id_router_002:sink_data
	wire         epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_rp_ready;                   // id_router_002:sink_ready -> epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent:rp_ready
	wire         uart_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                               // uart_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_003:sink_endofpacket
	wire         uart_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                                     // uart_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_003:sink_valid
	wire         uart_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                             // uart_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_003:sink_startofpacket
	wire  [93:0] uart_s1_translator_avalon_universal_slave_0_agent_rp_data;                                                      // uart_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_003:sink_data
	wire         uart_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                                     // id_router_003:sink_ready -> uart_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;                           // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_004:sink_endofpacket
	wire         jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid;                                 // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_004:sink_valid
	wire         jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;                         // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_004:sink_startofpacket
	wire  [93:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data;                                  // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_004:sink_data
	wire         jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready;                                 // id_router_004:sink_ready -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire         data_h_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                             // DATA_H_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_005:sink_endofpacket
	wire         data_h_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                                   // DATA_H_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_005:sink_valid
	wire         data_h_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                           // DATA_H_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_005:sink_startofpacket
	wire  [93:0] data_h_s1_translator_avalon_universal_slave_0_agent_rp_data;                                                    // DATA_H_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_005:sink_data
	wire         data_h_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                                   // id_router_005:sink_ready -> DATA_H_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                   // sysid_control_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_006:sink_endofpacket
	wire         sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_valid;                                         // sysid_control_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_006:sink_valid
	wire         sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                 // sysid_control_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_006:sink_startofpacket
	wire  [93:0] sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_data;                                          // sysid_control_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_006:sink_data
	wire         sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_ready;                                         // id_router_006:sink_ready -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire         data_l_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                             // DATA_L_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_007:sink_endofpacket
	wire         data_l_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                                   // DATA_L_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_007:sink_valid
	wire         data_l_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                           // DATA_L_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_007:sink_startofpacket
	wire  [93:0] data_l_s1_translator_avalon_universal_slave_0_agent_rp_data;                                                    // DATA_L_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_007:sink_data
	wire         data_l_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                                   // id_router_007:sink_ready -> DATA_L_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         pre_come_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                           // pre_come_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_008:sink_endofpacket
	wire         pre_come_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                                 // pre_come_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_008:sink_valid
	wire         pre_come_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                         // pre_come_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_008:sink_startofpacket
	wire  [93:0] pre_come_s1_translator_avalon_universal_slave_0_agent_rp_data;                                                  // pre_come_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_008:sink_data
	wire         pre_come_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                                 // id_router_008:sink_ready -> pre_come_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         tx_data_l_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                          // TX_DATA_L_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_009:sink_endofpacket
	wire         tx_data_l_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                                // TX_DATA_L_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_009:sink_valid
	wire         tx_data_l_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                        // TX_DATA_L_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_009:sink_startofpacket
	wire  [93:0] tx_data_l_s1_translator_avalon_universal_slave_0_agent_rp_data;                                                 // TX_DATA_L_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_009:sink_data
	wire         tx_data_l_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                                // id_router_009:sink_ready -> TX_DATA_L_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         tx_data_h_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                          // TX_DATA_H_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_010:sink_endofpacket
	wire         tx_data_h_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                                // TX_DATA_H_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_010:sink_valid
	wire         tx_data_h_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                        // TX_DATA_H_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_010:sink_startofpacket
	wire  [93:0] tx_data_h_s1_translator_avalon_universal_slave_0_agent_rp_data;                                                 // TX_DATA_H_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_010:sink_data
	wire         tx_data_h_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                                // id_router_010:sink_ready -> TX_DATA_H_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         tx_data_valid_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                      // TX_DATA_VALID_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_011:sink_endofpacket
	wire         tx_data_valid_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                            // TX_DATA_VALID_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_011:sink_valid
	wire         tx_data_valid_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                    // TX_DATA_VALID_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_011:sink_startofpacket
	wire  [93:0] tx_data_valid_s1_translator_avalon_universal_slave_0_agent_rp_data;                                             // TX_DATA_VALID_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_011:sink_data
	wire         tx_data_valid_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                            // id_router_011:sink_ready -> TX_DATA_VALID_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         addr_router_src_endofpacket;                                                                                    // addr_router:src_endofpacket -> limiter:cmd_sink_endofpacket
	wire         addr_router_src_valid;                                                                                          // addr_router:src_valid -> limiter:cmd_sink_valid
	wire         addr_router_src_startofpacket;                                                                                  // addr_router:src_startofpacket -> limiter:cmd_sink_startofpacket
	wire  [93:0] addr_router_src_data;                                                                                           // addr_router:src_data -> limiter:cmd_sink_data
	wire  [11:0] addr_router_src_channel;                                                                                        // addr_router:src_channel -> limiter:cmd_sink_channel
	wire         addr_router_src_ready;                                                                                          // limiter:cmd_sink_ready -> addr_router:src_ready
	wire         limiter_rsp_src_endofpacket;                                                                                    // limiter:rsp_src_endofpacket -> CPU_instruction_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire         limiter_rsp_src_valid;                                                                                          // limiter:rsp_src_valid -> CPU_instruction_master_translator_avalon_universal_master_0_agent:rp_valid
	wire         limiter_rsp_src_startofpacket;                                                                                  // limiter:rsp_src_startofpacket -> CPU_instruction_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [93:0] limiter_rsp_src_data;                                                                                           // limiter:rsp_src_data -> CPU_instruction_master_translator_avalon_universal_master_0_agent:rp_data
	wire  [11:0] limiter_rsp_src_channel;                                                                                        // limiter:rsp_src_channel -> CPU_instruction_master_translator_avalon_universal_master_0_agent:rp_channel
	wire         limiter_rsp_src_ready;                                                                                          // CPU_instruction_master_translator_avalon_universal_master_0_agent:rp_ready -> limiter:rsp_src_ready
	wire         addr_router_001_src_endofpacket;                                                                                // addr_router_001:src_endofpacket -> limiter_001:cmd_sink_endofpacket
	wire         addr_router_001_src_valid;                                                                                      // addr_router_001:src_valid -> limiter_001:cmd_sink_valid
	wire         addr_router_001_src_startofpacket;                                                                              // addr_router_001:src_startofpacket -> limiter_001:cmd_sink_startofpacket
	wire  [93:0] addr_router_001_src_data;                                                                                       // addr_router_001:src_data -> limiter_001:cmd_sink_data
	wire  [11:0] addr_router_001_src_channel;                                                                                    // addr_router_001:src_channel -> limiter_001:cmd_sink_channel
	wire         addr_router_001_src_ready;                                                                                      // limiter_001:cmd_sink_ready -> addr_router_001:src_ready
	wire         limiter_001_rsp_src_endofpacket;                                                                                // limiter_001:rsp_src_endofpacket -> CPU_data_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire         limiter_001_rsp_src_valid;                                                                                      // limiter_001:rsp_src_valid -> CPU_data_master_translator_avalon_universal_master_0_agent:rp_valid
	wire         limiter_001_rsp_src_startofpacket;                                                                              // limiter_001:rsp_src_startofpacket -> CPU_data_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [93:0] limiter_001_rsp_src_data;                                                                                       // limiter_001:rsp_src_data -> CPU_data_master_translator_avalon_universal_master_0_agent:rp_data
	wire  [11:0] limiter_001_rsp_src_channel;                                                                                    // limiter_001:rsp_src_channel -> CPU_data_master_translator_avalon_universal_master_0_agent:rp_channel
	wire         limiter_001_rsp_src_ready;                                                                                      // CPU_data_master_translator_avalon_universal_master_0_agent:rp_ready -> limiter_001:rsp_src_ready
	wire         rst_controller_reset_out_reset;                                                                                 // rst_controller:reset_out -> [CPU:reset_n, CPU_data_master_translator:reset, CPU_data_master_translator_avalon_universal_master_0_agent:reset, CPU_instruction_master_translator:reset, CPU_instruction_master_translator_avalon_universal_master_0_agent:reset, CPU_jtag_debug_module_translator:reset, CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:reset, CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, DATA_H:reset_n, DATA_H_s1_translator:reset, DATA_H_s1_translator_avalon_universal_slave_0_agent:reset, DATA_H_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, DATA_L:reset_n, DATA_L_s1_translator:reset, DATA_L_s1_translator_avalon_universal_slave_0_agent:reset, DATA_L_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, RAM:reset, RAM_s1_translator:reset, RAM_s1_translator_avalon_universal_slave_0_agent:reset, RAM_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, TX_DATA_H:reset_n, TX_DATA_H_s1_translator:reset, TX_DATA_H_s1_translator_avalon_universal_slave_0_agent:reset, TX_DATA_H_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, TX_DATA_L:reset_n, TX_DATA_L_s1_translator:reset, TX_DATA_L_s1_translator_avalon_universal_slave_0_agent:reset, TX_DATA_L_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, TX_DATA_VALID:reset_n, TX_DATA_VALID_s1_translator:reset, TX_DATA_VALID_s1_translator_avalon_universal_slave_0_agent:reset, TX_DATA_VALID_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, addr_router:reset, addr_router_001:reset, cmd_xbar_demux:reset, cmd_xbar_demux_001:reset, cmd_xbar_mux:reset, cmd_xbar_mux_001:reset, cmd_xbar_mux_002:reset, epcs_flash_controller_0:reset_n, epcs_flash_controller_0_epcs_control_port_translator:reset, epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent:reset, epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, id_router:reset, id_router_001:reset, id_router_002:reset, id_router_003:reset, id_router_004:reset, id_router_005:reset, id_router_006:reset, id_router_007:reset, id_router_008:reset, id_router_009:reset, id_router_010:reset, id_router_011:reset, irq_mapper:reset, jtag_uart:rst_n, jtag_uart_avalon_jtag_slave_translator:reset, jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:reset, jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, limiter:reset, limiter_001:reset, pre_come:reset_n, pre_come_s1_translator:reset, pre_come_s1_translator_avalon_universal_slave_0_agent:reset, pre_come_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, rsp_xbar_demux:reset, rsp_xbar_demux_001:reset, rsp_xbar_demux_002:reset, rsp_xbar_demux_003:reset, rsp_xbar_demux_004:reset, rsp_xbar_demux_005:reset, rsp_xbar_demux_006:reset, rsp_xbar_demux_007:reset, rsp_xbar_demux_008:reset, rsp_xbar_demux_009:reset, rsp_xbar_demux_010:reset, rsp_xbar_demux_011:reset, rsp_xbar_mux:reset, rsp_xbar_mux_001:reset, sysid:reset_n, sysid_control_slave_translator:reset, sysid_control_slave_translator_avalon_universal_slave_0_agent:reset, sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, uart:reset_n, uart_s1_translator:reset, uart_s1_translator_avalon_universal_slave_0_agent:reset, uart_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset]
	wire         cpu_jtag_debug_module_reset_reset;                                                                              // CPU:jtag_debug_module_resetrequest -> rst_controller:reset_in1
	wire         cmd_xbar_demux_src0_endofpacket;                                                                                // cmd_xbar_demux:src0_endofpacket -> cmd_xbar_mux:sink0_endofpacket
	wire         cmd_xbar_demux_src0_valid;                                                                                      // cmd_xbar_demux:src0_valid -> cmd_xbar_mux:sink0_valid
	wire         cmd_xbar_demux_src0_startofpacket;                                                                              // cmd_xbar_demux:src0_startofpacket -> cmd_xbar_mux:sink0_startofpacket
	wire  [93:0] cmd_xbar_demux_src0_data;                                                                                       // cmd_xbar_demux:src0_data -> cmd_xbar_mux:sink0_data
	wire  [11:0] cmd_xbar_demux_src0_channel;                                                                                    // cmd_xbar_demux:src0_channel -> cmd_xbar_mux:sink0_channel
	wire         cmd_xbar_demux_src0_ready;                                                                                      // cmd_xbar_mux:sink0_ready -> cmd_xbar_demux:src0_ready
	wire         cmd_xbar_demux_src1_endofpacket;                                                                                // cmd_xbar_demux:src1_endofpacket -> cmd_xbar_mux_001:sink0_endofpacket
	wire         cmd_xbar_demux_src1_valid;                                                                                      // cmd_xbar_demux:src1_valid -> cmd_xbar_mux_001:sink0_valid
	wire         cmd_xbar_demux_src1_startofpacket;                                                                              // cmd_xbar_demux:src1_startofpacket -> cmd_xbar_mux_001:sink0_startofpacket
	wire  [93:0] cmd_xbar_demux_src1_data;                                                                                       // cmd_xbar_demux:src1_data -> cmd_xbar_mux_001:sink0_data
	wire  [11:0] cmd_xbar_demux_src1_channel;                                                                                    // cmd_xbar_demux:src1_channel -> cmd_xbar_mux_001:sink0_channel
	wire         cmd_xbar_demux_src1_ready;                                                                                      // cmd_xbar_mux_001:sink0_ready -> cmd_xbar_demux:src1_ready
	wire         cmd_xbar_demux_src2_endofpacket;                                                                                // cmd_xbar_demux:src2_endofpacket -> cmd_xbar_mux_002:sink0_endofpacket
	wire         cmd_xbar_demux_src2_valid;                                                                                      // cmd_xbar_demux:src2_valid -> cmd_xbar_mux_002:sink0_valid
	wire         cmd_xbar_demux_src2_startofpacket;                                                                              // cmd_xbar_demux:src2_startofpacket -> cmd_xbar_mux_002:sink0_startofpacket
	wire  [93:0] cmd_xbar_demux_src2_data;                                                                                       // cmd_xbar_demux:src2_data -> cmd_xbar_mux_002:sink0_data
	wire  [11:0] cmd_xbar_demux_src2_channel;                                                                                    // cmd_xbar_demux:src2_channel -> cmd_xbar_mux_002:sink0_channel
	wire         cmd_xbar_demux_src2_ready;                                                                                      // cmd_xbar_mux_002:sink0_ready -> cmd_xbar_demux:src2_ready
	wire         cmd_xbar_demux_001_src0_endofpacket;                                                                            // cmd_xbar_demux_001:src0_endofpacket -> cmd_xbar_mux:sink1_endofpacket
	wire         cmd_xbar_demux_001_src0_valid;                                                                                  // cmd_xbar_demux_001:src0_valid -> cmd_xbar_mux:sink1_valid
	wire         cmd_xbar_demux_001_src0_startofpacket;                                                                          // cmd_xbar_demux_001:src0_startofpacket -> cmd_xbar_mux:sink1_startofpacket
	wire  [93:0] cmd_xbar_demux_001_src0_data;                                                                                   // cmd_xbar_demux_001:src0_data -> cmd_xbar_mux:sink1_data
	wire  [11:0] cmd_xbar_demux_001_src0_channel;                                                                                // cmd_xbar_demux_001:src0_channel -> cmd_xbar_mux:sink1_channel
	wire         cmd_xbar_demux_001_src0_ready;                                                                                  // cmd_xbar_mux:sink1_ready -> cmd_xbar_demux_001:src0_ready
	wire         cmd_xbar_demux_001_src1_endofpacket;                                                                            // cmd_xbar_demux_001:src1_endofpacket -> cmd_xbar_mux_001:sink1_endofpacket
	wire         cmd_xbar_demux_001_src1_valid;                                                                                  // cmd_xbar_demux_001:src1_valid -> cmd_xbar_mux_001:sink1_valid
	wire         cmd_xbar_demux_001_src1_startofpacket;                                                                          // cmd_xbar_demux_001:src1_startofpacket -> cmd_xbar_mux_001:sink1_startofpacket
	wire  [93:0] cmd_xbar_demux_001_src1_data;                                                                                   // cmd_xbar_demux_001:src1_data -> cmd_xbar_mux_001:sink1_data
	wire  [11:0] cmd_xbar_demux_001_src1_channel;                                                                                // cmd_xbar_demux_001:src1_channel -> cmd_xbar_mux_001:sink1_channel
	wire         cmd_xbar_demux_001_src1_ready;                                                                                  // cmd_xbar_mux_001:sink1_ready -> cmd_xbar_demux_001:src1_ready
	wire         cmd_xbar_demux_001_src2_endofpacket;                                                                            // cmd_xbar_demux_001:src2_endofpacket -> cmd_xbar_mux_002:sink1_endofpacket
	wire         cmd_xbar_demux_001_src2_valid;                                                                                  // cmd_xbar_demux_001:src2_valid -> cmd_xbar_mux_002:sink1_valid
	wire         cmd_xbar_demux_001_src2_startofpacket;                                                                          // cmd_xbar_demux_001:src2_startofpacket -> cmd_xbar_mux_002:sink1_startofpacket
	wire  [93:0] cmd_xbar_demux_001_src2_data;                                                                                   // cmd_xbar_demux_001:src2_data -> cmd_xbar_mux_002:sink1_data
	wire  [11:0] cmd_xbar_demux_001_src2_channel;                                                                                // cmd_xbar_demux_001:src2_channel -> cmd_xbar_mux_002:sink1_channel
	wire         cmd_xbar_demux_001_src2_ready;                                                                                  // cmd_xbar_mux_002:sink1_ready -> cmd_xbar_demux_001:src2_ready
	wire         cmd_xbar_demux_001_src3_endofpacket;                                                                            // cmd_xbar_demux_001:src3_endofpacket -> uart_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_001_src3_valid;                                                                                  // cmd_xbar_demux_001:src3_valid -> uart_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_001_src3_startofpacket;                                                                          // cmd_xbar_demux_001:src3_startofpacket -> uart_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [93:0] cmd_xbar_demux_001_src3_data;                                                                                   // cmd_xbar_demux_001:src3_data -> uart_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire  [11:0] cmd_xbar_demux_001_src3_channel;                                                                                // cmd_xbar_demux_001:src3_channel -> uart_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_001_src4_endofpacket;                                                                            // cmd_xbar_demux_001:src4_endofpacket -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_001_src4_valid;                                                                                  // cmd_xbar_demux_001:src4_valid -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_001_src4_startofpacket;                                                                          // cmd_xbar_demux_001:src4_startofpacket -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [93:0] cmd_xbar_demux_001_src4_data;                                                                                   // cmd_xbar_demux_001:src4_data -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire  [11:0] cmd_xbar_demux_001_src4_channel;                                                                                // cmd_xbar_demux_001:src4_channel -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_001_src5_endofpacket;                                                                            // cmd_xbar_demux_001:src5_endofpacket -> DATA_H_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_001_src5_valid;                                                                                  // cmd_xbar_demux_001:src5_valid -> DATA_H_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_001_src5_startofpacket;                                                                          // cmd_xbar_demux_001:src5_startofpacket -> DATA_H_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [93:0] cmd_xbar_demux_001_src5_data;                                                                                   // cmd_xbar_demux_001:src5_data -> DATA_H_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire  [11:0] cmd_xbar_demux_001_src5_channel;                                                                                // cmd_xbar_demux_001:src5_channel -> DATA_H_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_001_src6_endofpacket;                                                                            // cmd_xbar_demux_001:src6_endofpacket -> sysid_control_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_001_src6_valid;                                                                                  // cmd_xbar_demux_001:src6_valid -> sysid_control_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_001_src6_startofpacket;                                                                          // cmd_xbar_demux_001:src6_startofpacket -> sysid_control_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [93:0] cmd_xbar_demux_001_src6_data;                                                                                   // cmd_xbar_demux_001:src6_data -> sysid_control_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire  [11:0] cmd_xbar_demux_001_src6_channel;                                                                                // cmd_xbar_demux_001:src6_channel -> sysid_control_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_001_src7_endofpacket;                                                                            // cmd_xbar_demux_001:src7_endofpacket -> DATA_L_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_001_src7_valid;                                                                                  // cmd_xbar_demux_001:src7_valid -> DATA_L_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_001_src7_startofpacket;                                                                          // cmd_xbar_demux_001:src7_startofpacket -> DATA_L_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [93:0] cmd_xbar_demux_001_src7_data;                                                                                   // cmd_xbar_demux_001:src7_data -> DATA_L_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire  [11:0] cmd_xbar_demux_001_src7_channel;                                                                                // cmd_xbar_demux_001:src7_channel -> DATA_L_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_001_src8_endofpacket;                                                                            // cmd_xbar_demux_001:src8_endofpacket -> pre_come_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_001_src8_valid;                                                                                  // cmd_xbar_demux_001:src8_valid -> pre_come_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_001_src8_startofpacket;                                                                          // cmd_xbar_demux_001:src8_startofpacket -> pre_come_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [93:0] cmd_xbar_demux_001_src8_data;                                                                                   // cmd_xbar_demux_001:src8_data -> pre_come_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire  [11:0] cmd_xbar_demux_001_src8_channel;                                                                                // cmd_xbar_demux_001:src8_channel -> pre_come_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_001_src9_endofpacket;                                                                            // cmd_xbar_demux_001:src9_endofpacket -> TX_DATA_L_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_001_src9_valid;                                                                                  // cmd_xbar_demux_001:src9_valid -> TX_DATA_L_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_001_src9_startofpacket;                                                                          // cmd_xbar_demux_001:src9_startofpacket -> TX_DATA_L_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [93:0] cmd_xbar_demux_001_src9_data;                                                                                   // cmd_xbar_demux_001:src9_data -> TX_DATA_L_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire  [11:0] cmd_xbar_demux_001_src9_channel;                                                                                // cmd_xbar_demux_001:src9_channel -> TX_DATA_L_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_001_src10_endofpacket;                                                                           // cmd_xbar_demux_001:src10_endofpacket -> TX_DATA_H_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_001_src10_valid;                                                                                 // cmd_xbar_demux_001:src10_valid -> TX_DATA_H_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_001_src10_startofpacket;                                                                         // cmd_xbar_demux_001:src10_startofpacket -> TX_DATA_H_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [93:0] cmd_xbar_demux_001_src10_data;                                                                                  // cmd_xbar_demux_001:src10_data -> TX_DATA_H_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire  [11:0] cmd_xbar_demux_001_src10_channel;                                                                               // cmd_xbar_demux_001:src10_channel -> TX_DATA_H_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_001_src11_endofpacket;                                                                           // cmd_xbar_demux_001:src11_endofpacket -> TX_DATA_VALID_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_001_src11_valid;                                                                                 // cmd_xbar_demux_001:src11_valid -> TX_DATA_VALID_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_001_src11_startofpacket;                                                                         // cmd_xbar_demux_001:src11_startofpacket -> TX_DATA_VALID_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [93:0] cmd_xbar_demux_001_src11_data;                                                                                  // cmd_xbar_demux_001:src11_data -> TX_DATA_VALID_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire  [11:0] cmd_xbar_demux_001_src11_channel;                                                                               // cmd_xbar_demux_001:src11_channel -> TX_DATA_VALID_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         rsp_xbar_demux_src0_endofpacket;                                                                                // rsp_xbar_demux:src0_endofpacket -> rsp_xbar_mux:sink0_endofpacket
	wire         rsp_xbar_demux_src0_valid;                                                                                      // rsp_xbar_demux:src0_valid -> rsp_xbar_mux:sink0_valid
	wire         rsp_xbar_demux_src0_startofpacket;                                                                              // rsp_xbar_demux:src0_startofpacket -> rsp_xbar_mux:sink0_startofpacket
	wire  [93:0] rsp_xbar_demux_src0_data;                                                                                       // rsp_xbar_demux:src0_data -> rsp_xbar_mux:sink0_data
	wire  [11:0] rsp_xbar_demux_src0_channel;                                                                                    // rsp_xbar_demux:src0_channel -> rsp_xbar_mux:sink0_channel
	wire         rsp_xbar_demux_src0_ready;                                                                                      // rsp_xbar_mux:sink0_ready -> rsp_xbar_demux:src0_ready
	wire         rsp_xbar_demux_src1_endofpacket;                                                                                // rsp_xbar_demux:src1_endofpacket -> rsp_xbar_mux_001:sink0_endofpacket
	wire         rsp_xbar_demux_src1_valid;                                                                                      // rsp_xbar_demux:src1_valid -> rsp_xbar_mux_001:sink0_valid
	wire         rsp_xbar_demux_src1_startofpacket;                                                                              // rsp_xbar_demux:src1_startofpacket -> rsp_xbar_mux_001:sink0_startofpacket
	wire  [93:0] rsp_xbar_demux_src1_data;                                                                                       // rsp_xbar_demux:src1_data -> rsp_xbar_mux_001:sink0_data
	wire  [11:0] rsp_xbar_demux_src1_channel;                                                                                    // rsp_xbar_demux:src1_channel -> rsp_xbar_mux_001:sink0_channel
	wire         rsp_xbar_demux_src1_ready;                                                                                      // rsp_xbar_mux_001:sink0_ready -> rsp_xbar_demux:src1_ready
	wire         rsp_xbar_demux_001_src0_endofpacket;                                                                            // rsp_xbar_demux_001:src0_endofpacket -> rsp_xbar_mux:sink1_endofpacket
	wire         rsp_xbar_demux_001_src0_valid;                                                                                  // rsp_xbar_demux_001:src0_valid -> rsp_xbar_mux:sink1_valid
	wire         rsp_xbar_demux_001_src0_startofpacket;                                                                          // rsp_xbar_demux_001:src0_startofpacket -> rsp_xbar_mux:sink1_startofpacket
	wire  [93:0] rsp_xbar_demux_001_src0_data;                                                                                   // rsp_xbar_demux_001:src0_data -> rsp_xbar_mux:sink1_data
	wire  [11:0] rsp_xbar_demux_001_src0_channel;                                                                                // rsp_xbar_demux_001:src0_channel -> rsp_xbar_mux:sink1_channel
	wire         rsp_xbar_demux_001_src0_ready;                                                                                  // rsp_xbar_mux:sink1_ready -> rsp_xbar_demux_001:src0_ready
	wire         rsp_xbar_demux_001_src1_endofpacket;                                                                            // rsp_xbar_demux_001:src1_endofpacket -> rsp_xbar_mux_001:sink1_endofpacket
	wire         rsp_xbar_demux_001_src1_valid;                                                                                  // rsp_xbar_demux_001:src1_valid -> rsp_xbar_mux_001:sink1_valid
	wire         rsp_xbar_demux_001_src1_startofpacket;                                                                          // rsp_xbar_demux_001:src1_startofpacket -> rsp_xbar_mux_001:sink1_startofpacket
	wire  [93:0] rsp_xbar_demux_001_src1_data;                                                                                   // rsp_xbar_demux_001:src1_data -> rsp_xbar_mux_001:sink1_data
	wire  [11:0] rsp_xbar_demux_001_src1_channel;                                                                                // rsp_xbar_demux_001:src1_channel -> rsp_xbar_mux_001:sink1_channel
	wire         rsp_xbar_demux_001_src1_ready;                                                                                  // rsp_xbar_mux_001:sink1_ready -> rsp_xbar_demux_001:src1_ready
	wire         rsp_xbar_demux_002_src0_endofpacket;                                                                            // rsp_xbar_demux_002:src0_endofpacket -> rsp_xbar_mux:sink2_endofpacket
	wire         rsp_xbar_demux_002_src0_valid;                                                                                  // rsp_xbar_demux_002:src0_valid -> rsp_xbar_mux:sink2_valid
	wire         rsp_xbar_demux_002_src0_startofpacket;                                                                          // rsp_xbar_demux_002:src0_startofpacket -> rsp_xbar_mux:sink2_startofpacket
	wire  [93:0] rsp_xbar_demux_002_src0_data;                                                                                   // rsp_xbar_demux_002:src0_data -> rsp_xbar_mux:sink2_data
	wire  [11:0] rsp_xbar_demux_002_src0_channel;                                                                                // rsp_xbar_demux_002:src0_channel -> rsp_xbar_mux:sink2_channel
	wire         rsp_xbar_demux_002_src0_ready;                                                                                  // rsp_xbar_mux:sink2_ready -> rsp_xbar_demux_002:src0_ready
	wire         rsp_xbar_demux_002_src1_endofpacket;                                                                            // rsp_xbar_demux_002:src1_endofpacket -> rsp_xbar_mux_001:sink2_endofpacket
	wire         rsp_xbar_demux_002_src1_valid;                                                                                  // rsp_xbar_demux_002:src1_valid -> rsp_xbar_mux_001:sink2_valid
	wire         rsp_xbar_demux_002_src1_startofpacket;                                                                          // rsp_xbar_demux_002:src1_startofpacket -> rsp_xbar_mux_001:sink2_startofpacket
	wire  [93:0] rsp_xbar_demux_002_src1_data;                                                                                   // rsp_xbar_demux_002:src1_data -> rsp_xbar_mux_001:sink2_data
	wire  [11:0] rsp_xbar_demux_002_src1_channel;                                                                                // rsp_xbar_demux_002:src1_channel -> rsp_xbar_mux_001:sink2_channel
	wire         rsp_xbar_demux_002_src1_ready;                                                                                  // rsp_xbar_mux_001:sink2_ready -> rsp_xbar_demux_002:src1_ready
	wire         rsp_xbar_demux_003_src0_endofpacket;                                                                            // rsp_xbar_demux_003:src0_endofpacket -> rsp_xbar_mux_001:sink3_endofpacket
	wire         rsp_xbar_demux_003_src0_valid;                                                                                  // rsp_xbar_demux_003:src0_valid -> rsp_xbar_mux_001:sink3_valid
	wire         rsp_xbar_demux_003_src0_startofpacket;                                                                          // rsp_xbar_demux_003:src0_startofpacket -> rsp_xbar_mux_001:sink3_startofpacket
	wire  [93:0] rsp_xbar_demux_003_src0_data;                                                                                   // rsp_xbar_demux_003:src0_data -> rsp_xbar_mux_001:sink3_data
	wire  [11:0] rsp_xbar_demux_003_src0_channel;                                                                                // rsp_xbar_demux_003:src0_channel -> rsp_xbar_mux_001:sink3_channel
	wire         rsp_xbar_demux_003_src0_ready;                                                                                  // rsp_xbar_mux_001:sink3_ready -> rsp_xbar_demux_003:src0_ready
	wire         rsp_xbar_demux_004_src0_endofpacket;                                                                            // rsp_xbar_demux_004:src0_endofpacket -> rsp_xbar_mux_001:sink4_endofpacket
	wire         rsp_xbar_demux_004_src0_valid;                                                                                  // rsp_xbar_demux_004:src0_valid -> rsp_xbar_mux_001:sink4_valid
	wire         rsp_xbar_demux_004_src0_startofpacket;                                                                          // rsp_xbar_demux_004:src0_startofpacket -> rsp_xbar_mux_001:sink4_startofpacket
	wire  [93:0] rsp_xbar_demux_004_src0_data;                                                                                   // rsp_xbar_demux_004:src0_data -> rsp_xbar_mux_001:sink4_data
	wire  [11:0] rsp_xbar_demux_004_src0_channel;                                                                                // rsp_xbar_demux_004:src0_channel -> rsp_xbar_mux_001:sink4_channel
	wire         rsp_xbar_demux_004_src0_ready;                                                                                  // rsp_xbar_mux_001:sink4_ready -> rsp_xbar_demux_004:src0_ready
	wire         rsp_xbar_demux_005_src0_endofpacket;                                                                            // rsp_xbar_demux_005:src0_endofpacket -> rsp_xbar_mux_001:sink5_endofpacket
	wire         rsp_xbar_demux_005_src0_valid;                                                                                  // rsp_xbar_demux_005:src0_valid -> rsp_xbar_mux_001:sink5_valid
	wire         rsp_xbar_demux_005_src0_startofpacket;                                                                          // rsp_xbar_demux_005:src0_startofpacket -> rsp_xbar_mux_001:sink5_startofpacket
	wire  [93:0] rsp_xbar_demux_005_src0_data;                                                                                   // rsp_xbar_demux_005:src0_data -> rsp_xbar_mux_001:sink5_data
	wire  [11:0] rsp_xbar_demux_005_src0_channel;                                                                                // rsp_xbar_demux_005:src0_channel -> rsp_xbar_mux_001:sink5_channel
	wire         rsp_xbar_demux_005_src0_ready;                                                                                  // rsp_xbar_mux_001:sink5_ready -> rsp_xbar_demux_005:src0_ready
	wire         rsp_xbar_demux_006_src0_endofpacket;                                                                            // rsp_xbar_demux_006:src0_endofpacket -> rsp_xbar_mux_001:sink6_endofpacket
	wire         rsp_xbar_demux_006_src0_valid;                                                                                  // rsp_xbar_demux_006:src0_valid -> rsp_xbar_mux_001:sink6_valid
	wire         rsp_xbar_demux_006_src0_startofpacket;                                                                          // rsp_xbar_demux_006:src0_startofpacket -> rsp_xbar_mux_001:sink6_startofpacket
	wire  [93:0] rsp_xbar_demux_006_src0_data;                                                                                   // rsp_xbar_demux_006:src0_data -> rsp_xbar_mux_001:sink6_data
	wire  [11:0] rsp_xbar_demux_006_src0_channel;                                                                                // rsp_xbar_demux_006:src0_channel -> rsp_xbar_mux_001:sink6_channel
	wire         rsp_xbar_demux_006_src0_ready;                                                                                  // rsp_xbar_mux_001:sink6_ready -> rsp_xbar_demux_006:src0_ready
	wire         rsp_xbar_demux_007_src0_endofpacket;                                                                            // rsp_xbar_demux_007:src0_endofpacket -> rsp_xbar_mux_001:sink7_endofpacket
	wire         rsp_xbar_demux_007_src0_valid;                                                                                  // rsp_xbar_demux_007:src0_valid -> rsp_xbar_mux_001:sink7_valid
	wire         rsp_xbar_demux_007_src0_startofpacket;                                                                          // rsp_xbar_demux_007:src0_startofpacket -> rsp_xbar_mux_001:sink7_startofpacket
	wire  [93:0] rsp_xbar_demux_007_src0_data;                                                                                   // rsp_xbar_demux_007:src0_data -> rsp_xbar_mux_001:sink7_data
	wire  [11:0] rsp_xbar_demux_007_src0_channel;                                                                                // rsp_xbar_demux_007:src0_channel -> rsp_xbar_mux_001:sink7_channel
	wire         rsp_xbar_demux_007_src0_ready;                                                                                  // rsp_xbar_mux_001:sink7_ready -> rsp_xbar_demux_007:src0_ready
	wire         rsp_xbar_demux_008_src0_endofpacket;                                                                            // rsp_xbar_demux_008:src0_endofpacket -> rsp_xbar_mux_001:sink8_endofpacket
	wire         rsp_xbar_demux_008_src0_valid;                                                                                  // rsp_xbar_demux_008:src0_valid -> rsp_xbar_mux_001:sink8_valid
	wire         rsp_xbar_demux_008_src0_startofpacket;                                                                          // rsp_xbar_demux_008:src0_startofpacket -> rsp_xbar_mux_001:sink8_startofpacket
	wire  [93:0] rsp_xbar_demux_008_src0_data;                                                                                   // rsp_xbar_demux_008:src0_data -> rsp_xbar_mux_001:sink8_data
	wire  [11:0] rsp_xbar_demux_008_src0_channel;                                                                                // rsp_xbar_demux_008:src0_channel -> rsp_xbar_mux_001:sink8_channel
	wire         rsp_xbar_demux_008_src0_ready;                                                                                  // rsp_xbar_mux_001:sink8_ready -> rsp_xbar_demux_008:src0_ready
	wire         rsp_xbar_demux_009_src0_endofpacket;                                                                            // rsp_xbar_demux_009:src0_endofpacket -> rsp_xbar_mux_001:sink9_endofpacket
	wire         rsp_xbar_demux_009_src0_valid;                                                                                  // rsp_xbar_demux_009:src0_valid -> rsp_xbar_mux_001:sink9_valid
	wire         rsp_xbar_demux_009_src0_startofpacket;                                                                          // rsp_xbar_demux_009:src0_startofpacket -> rsp_xbar_mux_001:sink9_startofpacket
	wire  [93:0] rsp_xbar_demux_009_src0_data;                                                                                   // rsp_xbar_demux_009:src0_data -> rsp_xbar_mux_001:sink9_data
	wire  [11:0] rsp_xbar_demux_009_src0_channel;                                                                                // rsp_xbar_demux_009:src0_channel -> rsp_xbar_mux_001:sink9_channel
	wire         rsp_xbar_demux_009_src0_ready;                                                                                  // rsp_xbar_mux_001:sink9_ready -> rsp_xbar_demux_009:src0_ready
	wire         rsp_xbar_demux_010_src0_endofpacket;                                                                            // rsp_xbar_demux_010:src0_endofpacket -> rsp_xbar_mux_001:sink10_endofpacket
	wire         rsp_xbar_demux_010_src0_valid;                                                                                  // rsp_xbar_demux_010:src0_valid -> rsp_xbar_mux_001:sink10_valid
	wire         rsp_xbar_demux_010_src0_startofpacket;                                                                          // rsp_xbar_demux_010:src0_startofpacket -> rsp_xbar_mux_001:sink10_startofpacket
	wire  [93:0] rsp_xbar_demux_010_src0_data;                                                                                   // rsp_xbar_demux_010:src0_data -> rsp_xbar_mux_001:sink10_data
	wire  [11:0] rsp_xbar_demux_010_src0_channel;                                                                                // rsp_xbar_demux_010:src0_channel -> rsp_xbar_mux_001:sink10_channel
	wire         rsp_xbar_demux_010_src0_ready;                                                                                  // rsp_xbar_mux_001:sink10_ready -> rsp_xbar_demux_010:src0_ready
	wire         rsp_xbar_demux_011_src0_endofpacket;                                                                            // rsp_xbar_demux_011:src0_endofpacket -> rsp_xbar_mux_001:sink11_endofpacket
	wire         rsp_xbar_demux_011_src0_valid;                                                                                  // rsp_xbar_demux_011:src0_valid -> rsp_xbar_mux_001:sink11_valid
	wire         rsp_xbar_demux_011_src0_startofpacket;                                                                          // rsp_xbar_demux_011:src0_startofpacket -> rsp_xbar_mux_001:sink11_startofpacket
	wire  [93:0] rsp_xbar_demux_011_src0_data;                                                                                   // rsp_xbar_demux_011:src0_data -> rsp_xbar_mux_001:sink11_data
	wire  [11:0] rsp_xbar_demux_011_src0_channel;                                                                                // rsp_xbar_demux_011:src0_channel -> rsp_xbar_mux_001:sink11_channel
	wire         rsp_xbar_demux_011_src0_ready;                                                                                  // rsp_xbar_mux_001:sink11_ready -> rsp_xbar_demux_011:src0_ready
	wire         limiter_cmd_src_endofpacket;                                                                                    // limiter:cmd_src_endofpacket -> cmd_xbar_demux:sink_endofpacket
	wire         limiter_cmd_src_startofpacket;                                                                                  // limiter:cmd_src_startofpacket -> cmd_xbar_demux:sink_startofpacket
	wire  [93:0] limiter_cmd_src_data;                                                                                           // limiter:cmd_src_data -> cmd_xbar_demux:sink_data
	wire  [11:0] limiter_cmd_src_channel;                                                                                        // limiter:cmd_src_channel -> cmd_xbar_demux:sink_channel
	wire         limiter_cmd_src_ready;                                                                                          // cmd_xbar_demux:sink_ready -> limiter:cmd_src_ready
	wire         rsp_xbar_mux_src_endofpacket;                                                                                   // rsp_xbar_mux:src_endofpacket -> limiter:rsp_sink_endofpacket
	wire         rsp_xbar_mux_src_valid;                                                                                         // rsp_xbar_mux:src_valid -> limiter:rsp_sink_valid
	wire         rsp_xbar_mux_src_startofpacket;                                                                                 // rsp_xbar_mux:src_startofpacket -> limiter:rsp_sink_startofpacket
	wire  [93:0] rsp_xbar_mux_src_data;                                                                                          // rsp_xbar_mux:src_data -> limiter:rsp_sink_data
	wire  [11:0] rsp_xbar_mux_src_channel;                                                                                       // rsp_xbar_mux:src_channel -> limiter:rsp_sink_channel
	wire         rsp_xbar_mux_src_ready;                                                                                         // limiter:rsp_sink_ready -> rsp_xbar_mux:src_ready
	wire         limiter_001_cmd_src_endofpacket;                                                                                // limiter_001:cmd_src_endofpacket -> cmd_xbar_demux_001:sink_endofpacket
	wire         limiter_001_cmd_src_startofpacket;                                                                              // limiter_001:cmd_src_startofpacket -> cmd_xbar_demux_001:sink_startofpacket
	wire  [93:0] limiter_001_cmd_src_data;                                                                                       // limiter_001:cmd_src_data -> cmd_xbar_demux_001:sink_data
	wire  [11:0] limiter_001_cmd_src_channel;                                                                                    // limiter_001:cmd_src_channel -> cmd_xbar_demux_001:sink_channel
	wire         limiter_001_cmd_src_ready;                                                                                      // cmd_xbar_demux_001:sink_ready -> limiter_001:cmd_src_ready
	wire         rsp_xbar_mux_001_src_endofpacket;                                                                               // rsp_xbar_mux_001:src_endofpacket -> limiter_001:rsp_sink_endofpacket
	wire         rsp_xbar_mux_001_src_valid;                                                                                     // rsp_xbar_mux_001:src_valid -> limiter_001:rsp_sink_valid
	wire         rsp_xbar_mux_001_src_startofpacket;                                                                             // rsp_xbar_mux_001:src_startofpacket -> limiter_001:rsp_sink_startofpacket
	wire  [93:0] rsp_xbar_mux_001_src_data;                                                                                      // rsp_xbar_mux_001:src_data -> limiter_001:rsp_sink_data
	wire  [11:0] rsp_xbar_mux_001_src_channel;                                                                                   // rsp_xbar_mux_001:src_channel -> limiter_001:rsp_sink_channel
	wire         rsp_xbar_mux_001_src_ready;                                                                                     // limiter_001:rsp_sink_ready -> rsp_xbar_mux_001:src_ready
	wire         cmd_xbar_mux_src_endofpacket;                                                                                   // cmd_xbar_mux:src_endofpacket -> CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_mux_src_valid;                                                                                         // cmd_xbar_mux:src_valid -> CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_mux_src_startofpacket;                                                                                 // cmd_xbar_mux:src_startofpacket -> CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [93:0] cmd_xbar_mux_src_data;                                                                                          // cmd_xbar_mux:src_data -> CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_data
	wire  [11:0] cmd_xbar_mux_src_channel;                                                                                       // cmd_xbar_mux:src_channel -> CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_mux_src_ready;                                                                                         // CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux:src_ready
	wire         id_router_src_endofpacket;                                                                                      // id_router:src_endofpacket -> rsp_xbar_demux:sink_endofpacket
	wire         id_router_src_valid;                                                                                            // id_router:src_valid -> rsp_xbar_demux:sink_valid
	wire         id_router_src_startofpacket;                                                                                    // id_router:src_startofpacket -> rsp_xbar_demux:sink_startofpacket
	wire  [93:0] id_router_src_data;                                                                                             // id_router:src_data -> rsp_xbar_demux:sink_data
	wire  [11:0] id_router_src_channel;                                                                                          // id_router:src_channel -> rsp_xbar_demux:sink_channel
	wire         id_router_src_ready;                                                                                            // rsp_xbar_demux:sink_ready -> id_router:src_ready
	wire         cmd_xbar_mux_001_src_endofpacket;                                                                               // cmd_xbar_mux_001:src_endofpacket -> RAM_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_mux_001_src_valid;                                                                                     // cmd_xbar_mux_001:src_valid -> RAM_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_mux_001_src_startofpacket;                                                                             // cmd_xbar_mux_001:src_startofpacket -> RAM_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [93:0] cmd_xbar_mux_001_src_data;                                                                                      // cmd_xbar_mux_001:src_data -> RAM_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire  [11:0] cmd_xbar_mux_001_src_channel;                                                                                   // cmd_xbar_mux_001:src_channel -> RAM_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_mux_001_src_ready;                                                                                     // RAM_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_001:src_ready
	wire         id_router_001_src_endofpacket;                                                                                  // id_router_001:src_endofpacket -> rsp_xbar_demux_001:sink_endofpacket
	wire         id_router_001_src_valid;                                                                                        // id_router_001:src_valid -> rsp_xbar_demux_001:sink_valid
	wire         id_router_001_src_startofpacket;                                                                                // id_router_001:src_startofpacket -> rsp_xbar_demux_001:sink_startofpacket
	wire  [93:0] id_router_001_src_data;                                                                                         // id_router_001:src_data -> rsp_xbar_demux_001:sink_data
	wire  [11:0] id_router_001_src_channel;                                                                                      // id_router_001:src_channel -> rsp_xbar_demux_001:sink_channel
	wire         id_router_001_src_ready;                                                                                        // rsp_xbar_demux_001:sink_ready -> id_router_001:src_ready
	wire         cmd_xbar_mux_002_src_endofpacket;                                                                               // cmd_xbar_mux_002:src_endofpacket -> epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_mux_002_src_valid;                                                                                     // cmd_xbar_mux_002:src_valid -> epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_mux_002_src_startofpacket;                                                                             // cmd_xbar_mux_002:src_startofpacket -> epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [93:0] cmd_xbar_mux_002_src_data;                                                                                      // cmd_xbar_mux_002:src_data -> epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent:cp_data
	wire  [11:0] cmd_xbar_mux_002_src_channel;                                                                                   // cmd_xbar_mux_002:src_channel -> epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_mux_002_src_ready;                                                                                     // epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_002:src_ready
	wire         id_router_002_src_endofpacket;                                                                                  // id_router_002:src_endofpacket -> rsp_xbar_demux_002:sink_endofpacket
	wire         id_router_002_src_valid;                                                                                        // id_router_002:src_valid -> rsp_xbar_demux_002:sink_valid
	wire         id_router_002_src_startofpacket;                                                                                // id_router_002:src_startofpacket -> rsp_xbar_demux_002:sink_startofpacket
	wire  [93:0] id_router_002_src_data;                                                                                         // id_router_002:src_data -> rsp_xbar_demux_002:sink_data
	wire  [11:0] id_router_002_src_channel;                                                                                      // id_router_002:src_channel -> rsp_xbar_demux_002:sink_channel
	wire         id_router_002_src_ready;                                                                                        // rsp_xbar_demux_002:sink_ready -> id_router_002:src_ready
	wire         cmd_xbar_demux_001_src3_ready;                                                                                  // uart_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src3_ready
	wire         id_router_003_src_endofpacket;                                                                                  // id_router_003:src_endofpacket -> rsp_xbar_demux_003:sink_endofpacket
	wire         id_router_003_src_valid;                                                                                        // id_router_003:src_valid -> rsp_xbar_demux_003:sink_valid
	wire         id_router_003_src_startofpacket;                                                                                // id_router_003:src_startofpacket -> rsp_xbar_demux_003:sink_startofpacket
	wire  [93:0] id_router_003_src_data;                                                                                         // id_router_003:src_data -> rsp_xbar_demux_003:sink_data
	wire  [11:0] id_router_003_src_channel;                                                                                      // id_router_003:src_channel -> rsp_xbar_demux_003:sink_channel
	wire         id_router_003_src_ready;                                                                                        // rsp_xbar_demux_003:sink_ready -> id_router_003:src_ready
	wire         cmd_xbar_demux_001_src4_ready;                                                                                  // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src4_ready
	wire         id_router_004_src_endofpacket;                                                                                  // id_router_004:src_endofpacket -> rsp_xbar_demux_004:sink_endofpacket
	wire         id_router_004_src_valid;                                                                                        // id_router_004:src_valid -> rsp_xbar_demux_004:sink_valid
	wire         id_router_004_src_startofpacket;                                                                                // id_router_004:src_startofpacket -> rsp_xbar_demux_004:sink_startofpacket
	wire  [93:0] id_router_004_src_data;                                                                                         // id_router_004:src_data -> rsp_xbar_demux_004:sink_data
	wire  [11:0] id_router_004_src_channel;                                                                                      // id_router_004:src_channel -> rsp_xbar_demux_004:sink_channel
	wire         id_router_004_src_ready;                                                                                        // rsp_xbar_demux_004:sink_ready -> id_router_004:src_ready
	wire         cmd_xbar_demux_001_src5_ready;                                                                                  // DATA_H_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src5_ready
	wire         id_router_005_src_endofpacket;                                                                                  // id_router_005:src_endofpacket -> rsp_xbar_demux_005:sink_endofpacket
	wire         id_router_005_src_valid;                                                                                        // id_router_005:src_valid -> rsp_xbar_demux_005:sink_valid
	wire         id_router_005_src_startofpacket;                                                                                // id_router_005:src_startofpacket -> rsp_xbar_demux_005:sink_startofpacket
	wire  [93:0] id_router_005_src_data;                                                                                         // id_router_005:src_data -> rsp_xbar_demux_005:sink_data
	wire  [11:0] id_router_005_src_channel;                                                                                      // id_router_005:src_channel -> rsp_xbar_demux_005:sink_channel
	wire         id_router_005_src_ready;                                                                                        // rsp_xbar_demux_005:sink_ready -> id_router_005:src_ready
	wire         cmd_xbar_demux_001_src6_ready;                                                                                  // sysid_control_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src6_ready
	wire         id_router_006_src_endofpacket;                                                                                  // id_router_006:src_endofpacket -> rsp_xbar_demux_006:sink_endofpacket
	wire         id_router_006_src_valid;                                                                                        // id_router_006:src_valid -> rsp_xbar_demux_006:sink_valid
	wire         id_router_006_src_startofpacket;                                                                                // id_router_006:src_startofpacket -> rsp_xbar_demux_006:sink_startofpacket
	wire  [93:0] id_router_006_src_data;                                                                                         // id_router_006:src_data -> rsp_xbar_demux_006:sink_data
	wire  [11:0] id_router_006_src_channel;                                                                                      // id_router_006:src_channel -> rsp_xbar_demux_006:sink_channel
	wire         id_router_006_src_ready;                                                                                        // rsp_xbar_demux_006:sink_ready -> id_router_006:src_ready
	wire         cmd_xbar_demux_001_src7_ready;                                                                                  // DATA_L_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src7_ready
	wire         id_router_007_src_endofpacket;                                                                                  // id_router_007:src_endofpacket -> rsp_xbar_demux_007:sink_endofpacket
	wire         id_router_007_src_valid;                                                                                        // id_router_007:src_valid -> rsp_xbar_demux_007:sink_valid
	wire         id_router_007_src_startofpacket;                                                                                // id_router_007:src_startofpacket -> rsp_xbar_demux_007:sink_startofpacket
	wire  [93:0] id_router_007_src_data;                                                                                         // id_router_007:src_data -> rsp_xbar_demux_007:sink_data
	wire  [11:0] id_router_007_src_channel;                                                                                      // id_router_007:src_channel -> rsp_xbar_demux_007:sink_channel
	wire         id_router_007_src_ready;                                                                                        // rsp_xbar_demux_007:sink_ready -> id_router_007:src_ready
	wire         cmd_xbar_demux_001_src8_ready;                                                                                  // pre_come_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src8_ready
	wire         id_router_008_src_endofpacket;                                                                                  // id_router_008:src_endofpacket -> rsp_xbar_demux_008:sink_endofpacket
	wire         id_router_008_src_valid;                                                                                        // id_router_008:src_valid -> rsp_xbar_demux_008:sink_valid
	wire         id_router_008_src_startofpacket;                                                                                // id_router_008:src_startofpacket -> rsp_xbar_demux_008:sink_startofpacket
	wire  [93:0] id_router_008_src_data;                                                                                         // id_router_008:src_data -> rsp_xbar_demux_008:sink_data
	wire  [11:0] id_router_008_src_channel;                                                                                      // id_router_008:src_channel -> rsp_xbar_demux_008:sink_channel
	wire         id_router_008_src_ready;                                                                                        // rsp_xbar_demux_008:sink_ready -> id_router_008:src_ready
	wire         cmd_xbar_demux_001_src9_ready;                                                                                  // TX_DATA_L_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src9_ready
	wire         id_router_009_src_endofpacket;                                                                                  // id_router_009:src_endofpacket -> rsp_xbar_demux_009:sink_endofpacket
	wire         id_router_009_src_valid;                                                                                        // id_router_009:src_valid -> rsp_xbar_demux_009:sink_valid
	wire         id_router_009_src_startofpacket;                                                                                // id_router_009:src_startofpacket -> rsp_xbar_demux_009:sink_startofpacket
	wire  [93:0] id_router_009_src_data;                                                                                         // id_router_009:src_data -> rsp_xbar_demux_009:sink_data
	wire  [11:0] id_router_009_src_channel;                                                                                      // id_router_009:src_channel -> rsp_xbar_demux_009:sink_channel
	wire         id_router_009_src_ready;                                                                                        // rsp_xbar_demux_009:sink_ready -> id_router_009:src_ready
	wire         cmd_xbar_demux_001_src10_ready;                                                                                 // TX_DATA_H_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src10_ready
	wire         id_router_010_src_endofpacket;                                                                                  // id_router_010:src_endofpacket -> rsp_xbar_demux_010:sink_endofpacket
	wire         id_router_010_src_valid;                                                                                        // id_router_010:src_valid -> rsp_xbar_demux_010:sink_valid
	wire         id_router_010_src_startofpacket;                                                                                // id_router_010:src_startofpacket -> rsp_xbar_demux_010:sink_startofpacket
	wire  [93:0] id_router_010_src_data;                                                                                         // id_router_010:src_data -> rsp_xbar_demux_010:sink_data
	wire  [11:0] id_router_010_src_channel;                                                                                      // id_router_010:src_channel -> rsp_xbar_demux_010:sink_channel
	wire         id_router_010_src_ready;                                                                                        // rsp_xbar_demux_010:sink_ready -> id_router_010:src_ready
	wire         cmd_xbar_demux_001_src11_ready;                                                                                 // TX_DATA_VALID_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src11_ready
	wire         id_router_011_src_endofpacket;                                                                                  // id_router_011:src_endofpacket -> rsp_xbar_demux_011:sink_endofpacket
	wire         id_router_011_src_valid;                                                                                        // id_router_011:src_valid -> rsp_xbar_demux_011:sink_valid
	wire         id_router_011_src_startofpacket;                                                                                // id_router_011:src_startofpacket -> rsp_xbar_demux_011:sink_startofpacket
	wire  [93:0] id_router_011_src_data;                                                                                         // id_router_011:src_data -> rsp_xbar_demux_011:sink_data
	wire  [11:0] id_router_011_src_channel;                                                                                      // id_router_011:src_channel -> rsp_xbar_demux_011:sink_channel
	wire         id_router_011_src_ready;                                                                                        // rsp_xbar_demux_011:sink_ready -> id_router_011:src_ready
	wire  [11:0] limiter_cmd_valid_data;                                                                                         // limiter:cmd_src_valid -> cmd_xbar_demux:sink_valid
	wire  [11:0] limiter_001_cmd_valid_data;                                                                                     // limiter_001:cmd_src_valid -> cmd_xbar_demux_001:sink_valid
	wire         irq_mapper_receiver0_irq;                                                                                       // jtag_uart:av_irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                                                                       // uart:irq -> irq_mapper:receiver1_irq
	wire         irq_mapper_receiver2_irq;                                                                                       // epcs_flash_controller_0:irq -> irq_mapper:receiver2_irq
	wire         irq_mapper_receiver3_irq;                                                                                       // pre_come:irq -> irq_mapper:receiver3_irq
	wire  [31:0] cpu_d_irq_irq;                                                                                                  // irq_mapper:sender_irq -> CPU:d_irq

	NIOS2_CPU cpu (
		.clk                                   (clk_clk),                                                            //                       clk.clk
		.reset_n                               (~rst_controller_reset_out_reset),                                    //                   reset_n.reset_n
		.d_address                             (cpu_data_master_address),                                            //               data_master.address
		.d_byteenable                          (cpu_data_master_byteenable),                                         //                          .byteenable
		.d_read                                (cpu_data_master_read),                                               //                          .read
		.d_readdata                            (cpu_data_master_readdata),                                           //                          .readdata
		.d_waitrequest                         (cpu_data_master_waitrequest),                                        //                          .waitrequest
		.d_write                               (cpu_data_master_write),                                              //                          .write
		.d_writedata                           (cpu_data_master_writedata),                                          //                          .writedata
		.d_readdatavalid                       (cpu_data_master_readdatavalid),                                      //                          .readdatavalid
		.jtag_debug_module_debugaccess_to_roms (cpu_data_master_debugaccess),                                        //                          .debugaccess
		.i_address                             (cpu_instruction_master_address),                                     //        instruction_master.address
		.i_read                                (cpu_instruction_master_read),                                        //                          .read
		.i_readdata                            (cpu_instruction_master_readdata),                                    //                          .readdata
		.i_waitrequest                         (cpu_instruction_master_waitrequest),                                 //                          .waitrequest
		.i_readdatavalid                       (cpu_instruction_master_readdatavalid),                               //                          .readdatavalid
		.d_irq                                 (cpu_d_irq_irq),                                                      //                     d_irq.irq
		.jtag_debug_module_resetrequest        (cpu_jtag_debug_module_reset_reset),                                  //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (cpu_jtag_debug_module_translator_avalon_anti_slave_0_address),       //         jtag_debug_module.address
		.jtag_debug_module_begintransfer       (cpu_jtag_debug_module_translator_avalon_anti_slave_0_begintransfer), //                          .begintransfer
		.jtag_debug_module_byteenable          (cpu_jtag_debug_module_translator_avalon_anti_slave_0_byteenable),    //                          .byteenable
		.jtag_debug_module_debugaccess         (cpu_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess),   //                          .debugaccess
		.jtag_debug_module_readdata            (cpu_jtag_debug_module_translator_avalon_anti_slave_0_readdata),      //                          .readdata
		.jtag_debug_module_select              (cpu_jtag_debug_module_translator_avalon_anti_slave_0_chipselect),    //                          .chipselect
		.jtag_debug_module_write               (cpu_jtag_debug_module_translator_avalon_anti_slave_0_write),         //                          .write
		.jtag_debug_module_writedata           (cpu_jtag_debug_module_translator_avalon_anti_slave_0_writedata),     //                          .writedata
		.no_ci_readra                          ()                                                                    // custom_instruction_master.readra
	);

	NIOS2_RAM ram (
		.clk        (clk_clk),                                          //   clk1.clk
		.address    (ram_s1_translator_avalon_anti_slave_0_address),    //     s1.address
		.chipselect (ram_s1_translator_avalon_anti_slave_0_chipselect), //       .chipselect
		.clken      (ram_s1_translator_avalon_anti_slave_0_clken),      //       .clken
		.readdata   (ram_s1_translator_avalon_anti_slave_0_readdata),   //       .readdata
		.write      (ram_s1_translator_avalon_anti_slave_0_write),      //       .write
		.writedata  (ram_s1_translator_avalon_anti_slave_0_writedata),  //       .writedata
		.byteenable (ram_s1_translator_avalon_anti_slave_0_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset)                    // reset1.reset
	);

	NIOS2_jtag_uart jtag_uart (
		.clk            (clk_clk),                                                                //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                                        //             reset.reset_n
		.av_chipselect  (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_address),     //                  .address
		.av_read_n      (~jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_read),       //                  .read_n
		.av_readdata    (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata),    //                  .readdata
		.av_write_n     (~jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_write),      //                  .write_n
		.av_writedata   (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata),   //                  .writedata
		.av_waitrequest (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                                                //               irq.irq
	);

	NIOS2_uart uart (
		.clk           (clk_clk),                                              //                 clk.clk
		.reset_n       (~rst_controller_reset_out_reset),                      //               reset.reset_n
		.address       (uart_s1_translator_avalon_anti_slave_0_address),       //                  s1.address
		.begintransfer (uart_s1_translator_avalon_anti_slave_0_begintransfer), //                    .begintransfer
		.chipselect    (uart_s1_translator_avalon_anti_slave_0_chipselect),    //                    .chipselect
		.read_n        (~uart_s1_translator_avalon_anti_slave_0_read),         //                    .read_n
		.write_n       (~uart_s1_translator_avalon_anti_slave_0_write),        //                    .write_n
		.writedata     (uart_s1_translator_avalon_anti_slave_0_writedata),     //                    .writedata
		.readdata      (uart_s1_translator_avalon_anti_slave_0_readdata),      //                    .readdata
		.dataavailable (),                                                     //                    .dataavailable
		.readyfordata  (),                                                     //                    .readyfordata
		.rxd           (uart_external_connection_rxd),                         // external_connection.export
		.txd           (uart_external_connection_txd),                         //                    .export
		.irq           (irq_mapper_receiver1_irq)                              //                 irq.irq
	);

	NIOS2_DATA_H data_h (
		.clk      (clk_clk),                                           //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                   //               reset.reset_n
		.address  (data_h_s1_translator_avalon_anti_slave_0_address),  //                  s1.address
		.readdata (data_h_s1_translator_avalon_anti_slave_0_readdata), //                    .readdata
		.in_port  (data_external_connection_export)                    // external_connection.export
	);

	NIOS2_epcs_flash_controller_0 epcs_flash_controller_0 (
		.clk           (clk_clk),                                                                             //               clk.clk
		.reset_n       (~rst_controller_reset_out_reset),                                                     //             reset.reset_n
		.address       (epcs_flash_controller_0_epcs_control_port_translator_avalon_anti_slave_0_address),    // epcs_control_port.address
		.chipselect    (epcs_flash_controller_0_epcs_control_port_translator_avalon_anti_slave_0_chipselect), //                  .chipselect
		.dataavailable (),                                                                                    //                  .dataavailable
		.endofpacket   (),                                                                                    //                  .endofpacket
		.read_n        (~epcs_flash_controller_0_epcs_control_port_translator_avalon_anti_slave_0_read),      //                  .read_n
		.readdata      (epcs_flash_controller_0_epcs_control_port_translator_avalon_anti_slave_0_readdata),   //                  .readdata
		.readyfordata  (),                                                                                    //                  .readyfordata
		.write_n       (~epcs_flash_controller_0_epcs_control_port_translator_avalon_anti_slave_0_write),     //                  .write_n
		.writedata     (epcs_flash_controller_0_epcs_control_port_translator_avalon_anti_slave_0_writedata),  //                  .writedata
		.irq           (irq_mapper_receiver2_irq),                                                            //               irq.irq
		.dclk          (epcs_flash_controller_0_external_dclk),                                               //          external.export
		.sce           (epcs_flash_controller_0_external_sce),                                                //                  .export
		.sdo           (epcs_flash_controller_0_external_sdo),                                                //                  .export
		.data0         (epcs_flash_controller_0_external_data0)                                               //                  .export
	);

	NIOS2_sysid sysid (
		.clock    (clk_clk),                                                     //           clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                             //         reset.reset_n
		.readdata (sysid_control_slave_translator_avalon_anti_slave_0_readdata), // control_slave.readdata
		.address  (sysid_control_slave_translator_avalon_anti_slave_0_address)   //              .address
	);

	NIOS2_DATA_L data_l (
		.clk      (clk_clk),                                           //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                   //               reset.reset_n
		.address  (data_l_s1_translator_avalon_anti_slave_0_address),  //                  s1.address
		.readdata (data_l_s1_translator_avalon_anti_slave_0_readdata), //                    .readdata
		.in_port  (data_l_external_connection_export)                  // external_connection.export
	);

	NIOS2_pre_come pre_come (
		.clk        (clk_clk),                                               //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                       //               reset.reset_n
		.address    (pre_come_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~pre_come_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (pre_come_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (pre_come_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (pre_come_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.in_port    (pre_come_external_connection_export),                   // external_connection.export
		.irq        (irq_mapper_receiver3_irq)                               //                 irq.irq
	);

	NIOS2_TX_DATA_L tx_data_l (
		.clk        (clk_clk),                                                //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                        //               reset.reset_n
		.address    (tx_data_l_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~tx_data_l_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (tx_data_l_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (tx_data_l_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (tx_data_l_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.out_port   (tx_data_l_external_connection_export)                    // external_connection.export
	);

	NIOS2_TX_DATA_H tx_data_h (
		.clk        (clk_clk),                                                //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                        //               reset.reset_n
		.address    (tx_data_h_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~tx_data_h_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (tx_data_h_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (tx_data_h_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (tx_data_h_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.out_port   (tx_data_h_external_connection_export)                    // external_connection.export
	);

	NIOS2_TX_DATA_VALID tx_data_valid (
		.clk        (clk_clk),                                                    //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                            //               reset.reset_n
		.address    (tx_data_valid_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~tx_data_valid_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (tx_data_valid_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (tx_data_valid_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (tx_data_valid_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.out_port   (tx_data_valid_external_connection_export)                    // external_connection.export
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (19),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (19),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (0),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (1),
		.USE_WAITREQUEST             (1),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (1),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) cpu_instruction_master_translator (
		.clk                   (clk_clk),                                                                   //                       clk.clk
		.reset                 (rst_controller_reset_out_reset),                                            //                     reset.reset
		.uav_address           (cpu_instruction_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount        (cpu_instruction_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read              (cpu_instruction_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write             (cpu_instruction_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest       (cpu_instruction_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid     (cpu_instruction_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable        (cpu_instruction_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata          (cpu_instruction_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata         (cpu_instruction_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock              (cpu_instruction_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess       (cpu_instruction_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address            (cpu_instruction_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest        (cpu_instruction_master_waitrequest),                                        //                          .waitrequest
		.av_read               (cpu_instruction_master_read),                                               //                          .read
		.av_readdata           (cpu_instruction_master_readdata),                                           //                          .readdata
		.av_readdatavalid      (cpu_instruction_master_readdatavalid),                                      //                          .readdatavalid
		.av_burstcount         (1'b1),                                                                      //               (terminated)
		.av_byteenable         (4'b1111),                                                                   //               (terminated)
		.av_beginbursttransfer (1'b0),                                                                      //               (terminated)
		.av_begintransfer      (1'b0),                                                                      //               (terminated)
		.av_chipselect         (1'b0),                                                                      //               (terminated)
		.av_write              (1'b0),                                                                      //               (terminated)
		.av_writedata          (32'b00000000000000000000000000000000),                                      //               (terminated)
		.av_lock               (1'b0),                                                                      //               (terminated)
		.av_debugaccess        (1'b0),                                                                      //               (terminated)
		.uav_clken             (),                                                                          //               (terminated)
		.av_clken              (1'b1)                                                                       //               (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (19),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (19),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (1),
		.USE_WAITREQUEST             (1),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) cpu_data_master_translator (
		.clk                   (clk_clk),                                                            //                       clk.clk
		.reset                 (rst_controller_reset_out_reset),                                     //                     reset.reset
		.uav_address           (cpu_data_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount        (cpu_data_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read              (cpu_data_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write             (cpu_data_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest       (cpu_data_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid     (cpu_data_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable        (cpu_data_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata          (cpu_data_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata         (cpu_data_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock              (cpu_data_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess       (cpu_data_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address            (cpu_data_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest        (cpu_data_master_waitrequest),                                        //                          .waitrequest
		.av_byteenable         (cpu_data_master_byteenable),                                         //                          .byteenable
		.av_read               (cpu_data_master_read),                                               //                          .read
		.av_readdata           (cpu_data_master_readdata),                                           //                          .readdata
		.av_readdatavalid      (cpu_data_master_readdatavalid),                                      //                          .readdatavalid
		.av_write              (cpu_data_master_write),                                              //                          .write
		.av_writedata          (cpu_data_master_writedata),                                          //                          .writedata
		.av_debugaccess        (cpu_data_master_debugaccess),                                        //                          .debugaccess
		.av_burstcount         (1'b1),                                                               //               (terminated)
		.av_beginbursttransfer (1'b0),                                                               //               (terminated)
		.av_begintransfer      (1'b0),                                                               //               (terminated)
		.av_chipselect         (1'b0),                                                               //               (terminated)
		.av_lock               (1'b0),                                                               //               (terminated)
		.uav_clken             (),                                                                   //               (terminated)
		.av_clken              (1'b1)                                                                //               (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (9),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (19),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) cpu_jtag_debug_module_translator (
		.clk                   (clk_clk),                                                                          //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                                   //                    reset.reset
		.uav_address           (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (cpu_jtag_debug_module_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (cpu_jtag_debug_module_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (cpu_jtag_debug_module_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (cpu_jtag_debug_module_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_begintransfer      (cpu_jtag_debug_module_translator_avalon_anti_slave_0_begintransfer),               //                         .begintransfer
		.av_byteenable         (cpu_jtag_debug_module_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_chipselect         (cpu_jtag_debug_module_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_debugaccess        (cpu_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess),                 //                         .debugaccess
		.av_read               (),                                                                                 //              (terminated)
		.av_beginbursttransfer (),                                                                                 //              (terminated)
		.av_burstcount         (),                                                                                 //              (terminated)
		.av_readdatavalid      (1'b0),                                                                             //              (terminated)
		.av_waitrequest        (1'b0),                                                                             //              (terminated)
		.av_writebyteenable    (),                                                                                 //              (terminated)
		.av_lock               (),                                                                                 //              (terminated)
		.av_clken              (),                                                                                 //              (terminated)
		.uav_clken             (1'b0),                                                                             //              (terminated)
		.av_outputenable       ()                                                                                  //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (15),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (19),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) ram_s1_translator (
		.clk                   (clk_clk),                                                           //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                    //                    reset.reset
		.uav_address           (ram_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (ram_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (ram_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (ram_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (ram_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (ram_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (ram_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (ram_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (ram_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (ram_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (ram_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (ram_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (ram_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (ram_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (ram_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable         (ram_s1_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_chipselect         (ram_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_clken              (ram_s1_translator_avalon_anti_slave_0_clken),                       //                         .clken
		.av_read               (),                                                                  //              (terminated)
		.av_begintransfer      (),                                                                  //              (terminated)
		.av_beginbursttransfer (),                                                                  //              (terminated)
		.av_burstcount         (),                                                                  //              (terminated)
		.av_readdatavalid      (1'b0),                                                              //              (terminated)
		.av_waitrequest        (1'b0),                                                              //              (terminated)
		.av_writebyteenable    (),                                                                  //              (terminated)
		.av_lock               (),                                                                  //              (terminated)
		.uav_clken             (1'b0),                                                              //              (terminated)
		.av_debugaccess        (),                                                                  //              (terminated)
		.av_outputenable       ()                                                                   //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (9),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (19),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (1),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) epcs_flash_controller_0_epcs_control_port_translator (
		.clk                   (clk_clk),                                                                                              //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                                                       //                    reset.reset
		.uav_address           (epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (epcs_flash_controller_0_epcs_control_port_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (epcs_flash_controller_0_epcs_control_port_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (epcs_flash_controller_0_epcs_control_port_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (epcs_flash_controller_0_epcs_control_port_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (epcs_flash_controller_0_epcs_control_port_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect         (epcs_flash_controller_0_epcs_control_port_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer      (),                                                                                                     //              (terminated)
		.av_beginbursttransfer (),                                                                                                     //              (terminated)
		.av_burstcount         (),                                                                                                     //              (terminated)
		.av_byteenable         (),                                                                                                     //              (terminated)
		.av_readdatavalid      (1'b0),                                                                                                 //              (terminated)
		.av_waitrequest        (1'b0),                                                                                                 //              (terminated)
		.av_writebyteenable    (),                                                                                                     //              (terminated)
		.av_lock               (),                                                                                                     //              (terminated)
		.av_clken              (),                                                                                                     //              (terminated)
		.uav_clken             (1'b0),                                                                                                 //              (terminated)
		.av_debugaccess        (),                                                                                                     //              (terminated)
		.av_outputenable       ()                                                                                                      //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (16),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (19),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (1),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) uart_s1_translator (
		.clk                   (clk_clk),                                                            //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                     //                    reset.reset
		.uav_address           (uart_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (uart_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (uart_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (uart_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (uart_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (uart_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (uart_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (uart_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (uart_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (uart_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (uart_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (uart_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (uart_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (uart_s1_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (uart_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (uart_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_begintransfer      (uart_s1_translator_avalon_anti_slave_0_begintransfer),               //                         .begintransfer
		.av_chipselect         (uart_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_beginbursttransfer (),                                                                   //              (terminated)
		.av_burstcount         (),                                                                   //              (terminated)
		.av_byteenable         (),                                                                   //              (terminated)
		.av_readdatavalid      (1'b0),                                                               //              (terminated)
		.av_waitrequest        (1'b0),                                                               //              (terminated)
		.av_writebyteenable    (),                                                                   //              (terminated)
		.av_lock               (),                                                                   //              (terminated)
		.av_clken              (),                                                                   //              (terminated)
		.uav_clken             (1'b0),                                                               //              (terminated)
		.av_debugaccess        (),                                                                   //              (terminated)
		.av_outputenable       ()                                                                    //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (19),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) jtag_uart_avalon_jtag_slave_translator (
		.clk                   (clk_clk),                                                                                //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                                         //                    reset.reset
		.uav_address           (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_waitrequest        (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_chipselect         (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer      (),                                                                                       //              (terminated)
		.av_beginbursttransfer (),                                                                                       //              (terminated)
		.av_burstcount         (),                                                                                       //              (terminated)
		.av_byteenable         (),                                                                                       //              (terminated)
		.av_readdatavalid      (1'b0),                                                                                   //              (terminated)
		.av_writebyteenable    (),                                                                                       //              (terminated)
		.av_lock               (),                                                                                       //              (terminated)
		.av_clken              (),                                                                                       //              (terminated)
		.uav_clken             (1'b0),                                                                                   //              (terminated)
		.av_debugaccess        (),                                                                                       //              (terminated)
		.av_outputenable       ()                                                                                        //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (19),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) data_h_s1_translator (
		.clk                   (clk_clk),                                                              //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                       //                    reset.reset
		.uav_address           (data_h_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (data_h_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (data_h_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (data_h_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (data_h_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (data_h_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (data_h_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (data_h_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (data_h_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (data_h_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (data_h_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (data_h_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_readdata           (data_h_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_write              (),                                                                     //              (terminated)
		.av_read               (),                                                                     //              (terminated)
		.av_writedata          (),                                                                     //              (terminated)
		.av_begintransfer      (),                                                                     //              (terminated)
		.av_beginbursttransfer (),                                                                     //              (terminated)
		.av_burstcount         (),                                                                     //              (terminated)
		.av_byteenable         (),                                                                     //              (terminated)
		.av_readdatavalid      (1'b0),                                                                 //              (terminated)
		.av_waitrequest        (1'b0),                                                                 //              (terminated)
		.av_writebyteenable    (),                                                                     //              (terminated)
		.av_lock               (),                                                                     //              (terminated)
		.av_chipselect         (),                                                                     //              (terminated)
		.av_clken              (),                                                                     //              (terminated)
		.uav_clken             (1'b0),                                                                 //              (terminated)
		.av_debugaccess        (),                                                                     //              (terminated)
		.av_outputenable       ()                                                                      //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (19),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) sysid_control_slave_translator (
		.clk                   (clk_clk),                                                                        //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                                 //                    reset.reset
		.uav_address           (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (sysid_control_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_readdata           (sysid_control_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_write              (),                                                                               //              (terminated)
		.av_read               (),                                                                               //              (terminated)
		.av_writedata          (),                                                                               //              (terminated)
		.av_begintransfer      (),                                                                               //              (terminated)
		.av_beginbursttransfer (),                                                                               //              (terminated)
		.av_burstcount         (),                                                                               //              (terminated)
		.av_byteenable         (),                                                                               //              (terminated)
		.av_readdatavalid      (1'b0),                                                                           //              (terminated)
		.av_waitrequest        (1'b0),                                                                           //              (terminated)
		.av_writebyteenable    (),                                                                               //              (terminated)
		.av_lock               (),                                                                               //              (terminated)
		.av_chipselect         (),                                                                               //              (terminated)
		.av_clken              (),                                                                               //              (terminated)
		.uav_clken             (1'b0),                                                                           //              (terminated)
		.av_debugaccess        (),                                                                               //              (terminated)
		.av_outputenable       ()                                                                                //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (19),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) data_l_s1_translator (
		.clk                   (clk_clk),                                                              //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                       //                    reset.reset
		.uav_address           (data_l_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (data_l_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (data_l_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (data_l_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (data_l_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (data_l_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (data_l_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (data_l_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (data_l_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (data_l_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (data_l_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (data_l_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_readdata           (data_l_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_write              (),                                                                     //              (terminated)
		.av_read               (),                                                                     //              (terminated)
		.av_writedata          (),                                                                     //              (terminated)
		.av_begintransfer      (),                                                                     //              (terminated)
		.av_beginbursttransfer (),                                                                     //              (terminated)
		.av_burstcount         (),                                                                     //              (terminated)
		.av_byteenable         (),                                                                     //              (terminated)
		.av_readdatavalid      (1'b0),                                                                 //              (terminated)
		.av_waitrequest        (1'b0),                                                                 //              (terminated)
		.av_writebyteenable    (),                                                                     //              (terminated)
		.av_lock               (),                                                                     //              (terminated)
		.av_chipselect         (),                                                                     //              (terminated)
		.av_clken              (),                                                                     //              (terminated)
		.uav_clken             (1'b0),                                                                 //              (terminated)
		.av_debugaccess        (),                                                                     //              (terminated)
		.av_outputenable       ()                                                                      //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (19),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) pre_come_s1_translator (
		.clk                   (clk_clk),                                                                //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                         //                    reset.reset
		.uav_address           (pre_come_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (pre_come_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (pre_come_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (pre_come_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (pre_come_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (pre_come_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (pre_come_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (pre_come_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (pre_come_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (pre_come_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (pre_come_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (pre_come_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (pre_come_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (pre_come_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (pre_come_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect         (pre_come_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read               (),                                                                       //              (terminated)
		.av_begintransfer      (),                                                                       //              (terminated)
		.av_beginbursttransfer (),                                                                       //              (terminated)
		.av_burstcount         (),                                                                       //              (terminated)
		.av_byteenable         (),                                                                       //              (terminated)
		.av_readdatavalid      (1'b0),                                                                   //              (terminated)
		.av_waitrequest        (1'b0),                                                                   //              (terminated)
		.av_writebyteenable    (),                                                                       //              (terminated)
		.av_lock               (),                                                                       //              (terminated)
		.av_clken              (),                                                                       //              (terminated)
		.uav_clken             (1'b0),                                                                   //              (terminated)
		.av_debugaccess        (),                                                                       //              (terminated)
		.av_outputenable       ()                                                                        //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (19),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) tx_data_l_s1_translator (
		.clk                   (clk_clk),                                                                 //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                          //                    reset.reset
		.uav_address           (tx_data_l_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (tx_data_l_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (tx_data_l_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (tx_data_l_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (tx_data_l_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (tx_data_l_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (tx_data_l_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (tx_data_l_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (tx_data_l_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (tx_data_l_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (tx_data_l_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (tx_data_l_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (tx_data_l_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (tx_data_l_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (tx_data_l_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect         (tx_data_l_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read               (),                                                                        //              (terminated)
		.av_begintransfer      (),                                                                        //              (terminated)
		.av_beginbursttransfer (),                                                                        //              (terminated)
		.av_burstcount         (),                                                                        //              (terminated)
		.av_byteenable         (),                                                                        //              (terminated)
		.av_readdatavalid      (1'b0),                                                                    //              (terminated)
		.av_waitrequest        (1'b0),                                                                    //              (terminated)
		.av_writebyteenable    (),                                                                        //              (terminated)
		.av_lock               (),                                                                        //              (terminated)
		.av_clken              (),                                                                        //              (terminated)
		.uav_clken             (1'b0),                                                                    //              (terminated)
		.av_debugaccess        (),                                                                        //              (terminated)
		.av_outputenable       ()                                                                         //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (19),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) tx_data_h_s1_translator (
		.clk                   (clk_clk),                                                                 //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                          //                    reset.reset
		.uav_address           (tx_data_h_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (tx_data_h_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (tx_data_h_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (tx_data_h_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (tx_data_h_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (tx_data_h_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (tx_data_h_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (tx_data_h_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (tx_data_h_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (tx_data_h_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (tx_data_h_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (tx_data_h_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (tx_data_h_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (tx_data_h_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (tx_data_h_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect         (tx_data_h_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read               (),                                                                        //              (terminated)
		.av_begintransfer      (),                                                                        //              (terminated)
		.av_beginbursttransfer (),                                                                        //              (terminated)
		.av_burstcount         (),                                                                        //              (terminated)
		.av_byteenable         (),                                                                        //              (terminated)
		.av_readdatavalid      (1'b0),                                                                    //              (terminated)
		.av_waitrequest        (1'b0),                                                                    //              (terminated)
		.av_writebyteenable    (),                                                                        //              (terminated)
		.av_lock               (),                                                                        //              (terminated)
		.av_clken              (),                                                                        //              (terminated)
		.uav_clken             (1'b0),                                                                    //              (terminated)
		.av_debugaccess        (),                                                                        //              (terminated)
		.av_outputenable       ()                                                                         //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (19),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) tx_data_valid_s1_translator (
		.clk                   (clk_clk),                                                                     //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                              //                    reset.reset
		.uav_address           (tx_data_valid_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (tx_data_valid_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (tx_data_valid_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (tx_data_valid_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (tx_data_valid_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (tx_data_valid_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (tx_data_valid_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (tx_data_valid_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (tx_data_valid_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (tx_data_valid_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (tx_data_valid_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (tx_data_valid_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (tx_data_valid_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (tx_data_valid_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (tx_data_valid_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect         (tx_data_valid_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read               (),                                                                            //              (terminated)
		.av_begintransfer      (),                                                                            //              (terminated)
		.av_beginbursttransfer (),                                                                            //              (terminated)
		.av_burstcount         (),                                                                            //              (terminated)
		.av_byteenable         (),                                                                            //              (terminated)
		.av_readdatavalid      (1'b0),                                                                        //              (terminated)
		.av_waitrequest        (1'b0),                                                                        //              (terminated)
		.av_writebyteenable    (),                                                                            //              (terminated)
		.av_lock               (),                                                                            //              (terminated)
		.av_clken              (),                                                                            //              (terminated)
		.uav_clken             (1'b0),                                                                        //              (terminated)
		.av_debugaccess        (),                                                                            //              (terminated)
		.av_outputenable       ()                                                                             //              (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (87),
		.PKT_PROTECTION_L          (85),
		.PKT_BEGIN_BURST           (74),
		.PKT_BURSTWRAP_H           (66),
		.PKT_BURSTWRAP_L           (64),
		.PKT_BURST_SIZE_H          (69),
		.PKT_BURST_SIZE_L          (67),
		.PKT_BURST_TYPE_H          (71),
		.PKT_BURST_TYPE_L          (70),
		.PKT_BYTE_CNT_H            (63),
		.PKT_BYTE_CNT_L            (61),
		.PKT_ADDR_H                (54),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (55),
		.PKT_TRANS_POSTED          (56),
		.PKT_TRANS_WRITE           (57),
		.PKT_TRANS_READ            (58),
		.PKT_TRANS_LOCK            (59),
		.PKT_TRANS_EXCLUSIVE       (60),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (79),
		.PKT_SRC_ID_L              (76),
		.PKT_DEST_ID_H             (83),
		.PKT_DEST_ID_L             (80),
		.PKT_THREAD_ID_H           (84),
		.PKT_THREAD_ID_L           (84),
		.PKT_CACHE_H               (91),
		.PKT_CACHE_L               (88),
		.PKT_DATA_SIDEBAND_H       (73),
		.PKT_DATA_SIDEBAND_L       (73),
		.PKT_QOS_H                 (75),
		.PKT_QOS_L                 (75),
		.PKT_ADDR_SIDEBAND_H       (72),
		.PKT_ADDR_SIDEBAND_L       (72),
		.ST_DATA_W                 (94),
		.ST_CHANNEL_W              (12),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (0),
		.BURSTWRAP_VALUE           (3),
		.CACHE_VALUE               (4'b0000)
	) cpu_instruction_master_translator_avalon_universal_master_0_agent (
		.clk              (clk_clk),                                                                            //       clk.clk
		.reset            (rst_controller_reset_out_reset),                                                     // clk_reset.reset
		.av_address       (cpu_instruction_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write         (cpu_instruction_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read          (cpu_instruction_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata     (cpu_instruction_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata      (cpu_instruction_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest   (cpu_instruction_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid (cpu_instruction_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable    (cpu_instruction_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount    (cpu_instruction_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess   (cpu_instruction_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock          (cpu_instruction_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid         (cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data          (cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket (cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket   (cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready         (cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid         (limiter_rsp_src_valid),                                                              //        rp.valid
		.rp_data          (limiter_rsp_src_data),                                                               //          .data
		.rp_channel       (limiter_rsp_src_channel),                                                            //          .channel
		.rp_startofpacket (limiter_rsp_src_startofpacket),                                                      //          .startofpacket
		.rp_endofpacket   (limiter_rsp_src_endofpacket),                                                        //          .endofpacket
		.rp_ready         (limiter_rsp_src_ready)                                                               //          .ready
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (87),
		.PKT_PROTECTION_L          (85),
		.PKT_BEGIN_BURST           (74),
		.PKT_BURSTWRAP_H           (66),
		.PKT_BURSTWRAP_L           (64),
		.PKT_BURST_SIZE_H          (69),
		.PKT_BURST_SIZE_L          (67),
		.PKT_BURST_TYPE_H          (71),
		.PKT_BURST_TYPE_L          (70),
		.PKT_BYTE_CNT_H            (63),
		.PKT_BYTE_CNT_L            (61),
		.PKT_ADDR_H                (54),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (55),
		.PKT_TRANS_POSTED          (56),
		.PKT_TRANS_WRITE           (57),
		.PKT_TRANS_READ            (58),
		.PKT_TRANS_LOCK            (59),
		.PKT_TRANS_EXCLUSIVE       (60),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (79),
		.PKT_SRC_ID_L              (76),
		.PKT_DEST_ID_H             (83),
		.PKT_DEST_ID_L             (80),
		.PKT_THREAD_ID_H           (84),
		.PKT_THREAD_ID_L           (84),
		.PKT_CACHE_H               (91),
		.PKT_CACHE_L               (88),
		.PKT_DATA_SIDEBAND_H       (73),
		.PKT_DATA_SIDEBAND_L       (73),
		.PKT_QOS_H                 (75),
		.PKT_QOS_L                 (75),
		.PKT_ADDR_SIDEBAND_H       (72),
		.PKT_ADDR_SIDEBAND_L       (72),
		.ST_DATA_W                 (94),
		.ST_CHANNEL_W              (12),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (1),
		.BURSTWRAP_VALUE           (7),
		.CACHE_VALUE               (4'b0000)
	) cpu_data_master_translator_avalon_universal_master_0_agent (
		.clk              (clk_clk),                                                                     //       clk.clk
		.reset            (rst_controller_reset_out_reset),                                              // clk_reset.reset
		.av_address       (cpu_data_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write         (cpu_data_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read          (cpu_data_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata     (cpu_data_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata      (cpu_data_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest   (cpu_data_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid (cpu_data_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable    (cpu_data_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount    (cpu_data_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess   (cpu_data_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock          (cpu_data_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid         (cpu_data_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data          (cpu_data_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket (cpu_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket   (cpu_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready         (cpu_data_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid         (limiter_001_rsp_src_valid),                                                   //        rp.valid
		.rp_data          (limiter_001_rsp_src_data),                                                    //          .data
		.rp_channel       (limiter_001_rsp_src_channel),                                                 //          .channel
		.rp_startofpacket (limiter_001_rsp_src_startofpacket),                                           //          .startofpacket
		.rp_endofpacket   (limiter_001_rsp_src_endofpacket),                                             //          .endofpacket
		.rp_ready         (limiter_001_rsp_src_ready)                                                    //          .ready
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (74),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (54),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (55),
		.PKT_TRANS_POSTED          (56),
		.PKT_TRANS_WRITE           (57),
		.PKT_TRANS_READ            (58),
		.PKT_TRANS_LOCK            (59),
		.PKT_SRC_ID_H              (79),
		.PKT_SRC_ID_L              (76),
		.PKT_DEST_ID_H             (83),
		.PKT_DEST_ID_L             (80),
		.PKT_BURSTWRAP_H           (66),
		.PKT_BURSTWRAP_L           (64),
		.PKT_BYTE_CNT_H            (63),
		.PKT_BYTE_CNT_L            (61),
		.PKT_PROTECTION_H          (87),
		.PKT_PROTECTION_L          (85),
		.PKT_RESPONSE_STATUS_H     (93),
		.PKT_RESPONSE_STATUS_L     (92),
		.PKT_BURST_SIZE_H          (69),
		.PKT_BURST_SIZE_L          (67),
		.ST_CHANNEL_W              (12),
		.ST_DATA_W                 (94),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                    //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                             //       clk_reset.reset
		.m0_address              (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_src_ready),                                                                     //              cp.ready
		.cp_valid                (cmd_xbar_mux_src_valid),                                                                     //                .valid
		.cp_data                 (cmd_xbar_mux_src_data),                                                                      //                .data
		.cp_startofpacket        (cmd_xbar_mux_src_startofpacket),                                                             //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_src_endofpacket),                                                               //                .endofpacket
		.cp_channel              (cmd_xbar_mux_src_channel),                                                                   //                .channel
		.rf_sink_ready           (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (95),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                    //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                             // clk_reset.reset
		.in_data           (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                      // (terminated)
		.csr_read          (1'b0),                                                                                       // (terminated)
		.csr_write         (1'b0),                                                                                       // (terminated)
		.csr_readdata      (),                                                                                           // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                       // (terminated)
		.almost_full_data  (),                                                                                           // (terminated)
		.almost_empty_data (),                                                                                           // (terminated)
		.in_empty          (1'b0),                                                                                       // (terminated)
		.out_empty         (),                                                                                           // (terminated)
		.in_error          (1'b0),                                                                                       // (terminated)
		.out_error         (),                                                                                           // (terminated)
		.in_channel        (1'b0),                                                                                       // (terminated)
		.out_channel       ()                                                                                            // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (74),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (54),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (55),
		.PKT_TRANS_POSTED          (56),
		.PKT_TRANS_WRITE           (57),
		.PKT_TRANS_READ            (58),
		.PKT_TRANS_LOCK            (59),
		.PKT_SRC_ID_H              (79),
		.PKT_SRC_ID_L              (76),
		.PKT_DEST_ID_H             (83),
		.PKT_DEST_ID_L             (80),
		.PKT_BURSTWRAP_H           (66),
		.PKT_BURSTWRAP_L           (64),
		.PKT_BYTE_CNT_H            (63),
		.PKT_BYTE_CNT_L            (61),
		.PKT_PROTECTION_H          (87),
		.PKT_PROTECTION_L          (85),
		.PKT_RESPONSE_STATUS_H     (93),
		.PKT_RESPONSE_STATUS_L     (92),
		.PKT_BURST_SIZE_H          (69),
		.PKT_BURST_SIZE_L          (67),
		.ST_CHANNEL_W              (12),
		.ST_DATA_W                 (94),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) ram_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                     //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                              //       clk_reset.reset
		.m0_address              (ram_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (ram_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (ram_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (ram_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (ram_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (ram_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (ram_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (ram_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (ram_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (ram_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (ram_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (ram_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (ram_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (ram_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (ram_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (ram_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_001_src_ready),                                                  //              cp.ready
		.cp_valid                (cmd_xbar_mux_001_src_valid),                                                  //                .valid
		.cp_data                 (cmd_xbar_mux_001_src_data),                                                   //                .data
		.cp_startofpacket        (cmd_xbar_mux_001_src_startofpacket),                                          //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_001_src_endofpacket),                                            //                .endofpacket
		.cp_channel              (cmd_xbar_mux_001_src_channel),                                                //                .channel
		.rf_sink_ready           (ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (ram_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (ram_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (ram_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (ram_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (ram_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (ram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (ram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (ram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (ram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (ram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (ram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (95),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                     //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                              // clk_reset.reset
		.in_data           (ram_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (ram_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (ram_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (ram_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (ram_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                       // (terminated)
		.csr_read          (1'b0),                                                                        // (terminated)
		.csr_write         (1'b0),                                                                        // (terminated)
		.csr_readdata      (),                                                                            // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                        // (terminated)
		.almost_full_data  (),                                                                            // (terminated)
		.almost_empty_data (),                                                                            // (terminated)
		.in_empty          (1'b0),                                                                        // (terminated)
		.out_empty         (),                                                                            // (terminated)
		.in_error          (1'b0),                                                                        // (terminated)
		.out_error         (),                                                                            // (terminated)
		.in_channel        (1'b0),                                                                        // (terminated)
		.out_channel       ()                                                                             // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (74),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (54),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (55),
		.PKT_TRANS_POSTED          (56),
		.PKT_TRANS_WRITE           (57),
		.PKT_TRANS_READ            (58),
		.PKT_TRANS_LOCK            (59),
		.PKT_SRC_ID_H              (79),
		.PKT_SRC_ID_L              (76),
		.PKT_DEST_ID_H             (83),
		.PKT_DEST_ID_L             (80),
		.PKT_BURSTWRAP_H           (66),
		.PKT_BURSTWRAP_L           (64),
		.PKT_BYTE_CNT_H            (63),
		.PKT_BYTE_CNT_L            (61),
		.PKT_PROTECTION_H          (87),
		.PKT_PROTECTION_L          (85),
		.PKT_RESPONSE_STATUS_H     (93),
		.PKT_RESPONSE_STATUS_L     (92),
		.PKT_BURST_SIZE_H          (69),
		.PKT_BURST_SIZE_L          (67),
		.ST_CHANNEL_W              (12),
		.ST_DATA_W                 (94),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                                        //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                                                 //       clk_reset.reset
		.m0_address              (epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_002_src_ready),                                                                                     //              cp.ready
		.cp_valid                (cmd_xbar_mux_002_src_valid),                                                                                     //                .valid
		.cp_data                 (cmd_xbar_mux_002_src_data),                                                                                      //                .data
		.cp_startofpacket        (cmd_xbar_mux_002_src_startofpacket),                                                                             //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_002_src_endofpacket),                                                                               //                .endofpacket
		.cp_channel              (cmd_xbar_mux_002_src_channel),                                                                                   //                .channel
		.rf_sink_ready           (epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (95),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                                        //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                                                 // clk_reset.reset
		.in_data           (epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                                          // (terminated)
		.csr_read          (1'b0),                                                                                                           // (terminated)
		.csr_write         (1'b0),                                                                                                           // (terminated)
		.csr_readdata      (),                                                                                                               // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                                           // (terminated)
		.almost_full_data  (),                                                                                                               // (terminated)
		.almost_empty_data (),                                                                                                               // (terminated)
		.in_empty          (1'b0),                                                                                                           // (terminated)
		.out_empty         (),                                                                                                               // (terminated)
		.in_error          (1'b0),                                                                                                           // (terminated)
		.out_error         (),                                                                                                               // (terminated)
		.in_channel        (1'b0),                                                                                                           // (terminated)
		.out_channel       ()                                                                                                                // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (74),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (54),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (55),
		.PKT_TRANS_POSTED          (56),
		.PKT_TRANS_WRITE           (57),
		.PKT_TRANS_READ            (58),
		.PKT_TRANS_LOCK            (59),
		.PKT_SRC_ID_H              (79),
		.PKT_SRC_ID_L              (76),
		.PKT_DEST_ID_H             (83),
		.PKT_DEST_ID_L             (80),
		.PKT_BURSTWRAP_H           (66),
		.PKT_BURSTWRAP_L           (64),
		.PKT_BYTE_CNT_H            (63),
		.PKT_BYTE_CNT_L            (61),
		.PKT_PROTECTION_H          (87),
		.PKT_PROTECTION_L          (85),
		.PKT_RESPONSE_STATUS_H     (93),
		.PKT_RESPONSE_STATUS_L     (92),
		.PKT_BURST_SIZE_H          (69),
		.PKT_BURST_SIZE_L          (67),
		.ST_CHANNEL_W              (12),
		.ST_DATA_W                 (94),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) uart_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                      //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                               //       clk_reset.reset
		.m0_address              (uart_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (uart_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (uart_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (uart_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (uart_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (uart_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (uart_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (uart_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (uart_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (uart_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (uart_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (uart_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (uart_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (uart_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (uart_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (uart_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src3_ready),                                                //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src3_valid),                                                //                .valid
		.cp_data                 (cmd_xbar_demux_001_src3_data),                                                 //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src3_startofpacket),                                        //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src3_endofpacket),                                          //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src3_channel),                                              //                .channel
		.rf_sink_ready           (uart_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (uart_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (uart_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (uart_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (uart_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (uart_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (uart_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (uart_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (uart_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (uart_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (uart_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (uart_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (uart_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (uart_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (uart_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (uart_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (95),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) uart_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                      //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                               // clk_reset.reset
		.in_data           (uart_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (uart_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (uart_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (uart_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (uart_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (uart_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (uart_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (uart_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (uart_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (uart_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                        // (terminated)
		.csr_read          (1'b0),                                                                         // (terminated)
		.csr_write         (1'b0),                                                                         // (terminated)
		.csr_readdata      (),                                                                             // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                         // (terminated)
		.almost_full_data  (),                                                                             // (terminated)
		.almost_empty_data (),                                                                             // (terminated)
		.in_empty          (1'b0),                                                                         // (terminated)
		.out_empty         (),                                                                             // (terminated)
		.in_error          (1'b0),                                                                         // (terminated)
		.out_error         (),                                                                             // (terminated)
		.in_channel        (1'b0),                                                                         // (terminated)
		.out_channel       ()                                                                              // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (74),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (54),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (55),
		.PKT_TRANS_POSTED          (56),
		.PKT_TRANS_WRITE           (57),
		.PKT_TRANS_READ            (58),
		.PKT_TRANS_LOCK            (59),
		.PKT_SRC_ID_H              (79),
		.PKT_SRC_ID_L              (76),
		.PKT_DEST_ID_H             (83),
		.PKT_DEST_ID_L             (80),
		.PKT_BURSTWRAP_H           (66),
		.PKT_BURSTWRAP_L           (64),
		.PKT_BYTE_CNT_H            (63),
		.PKT_BYTE_CNT_L            (61),
		.PKT_PROTECTION_H          (87),
		.PKT_PROTECTION_L          (85),
		.PKT_RESPONSE_STATUS_H     (93),
		.PKT_RESPONSE_STATUS_L     (92),
		.PKT_BURST_SIZE_H          (69),
		.PKT_BURST_SIZE_L          (67),
		.ST_CHANNEL_W              (12),
		.ST_DATA_W                 (94),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                          //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                                   //       clk_reset.reset
		.m0_address              (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src4_ready),                                                                    //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src4_valid),                                                                    //                .valid
		.cp_data                 (cmd_xbar_demux_001_src4_data),                                                                     //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src4_startofpacket),                                                            //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src4_endofpacket),                                                              //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src4_channel),                                                                  //                .channel
		.rf_sink_ready           (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (95),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                          //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                                   // clk_reset.reset
		.in_data           (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                            // (terminated)
		.csr_read          (1'b0),                                                                                             // (terminated)
		.csr_write         (1'b0),                                                                                             // (terminated)
		.csr_readdata      (),                                                                                                 // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                             // (terminated)
		.almost_full_data  (),                                                                                                 // (terminated)
		.almost_empty_data (),                                                                                                 // (terminated)
		.in_empty          (1'b0),                                                                                             // (terminated)
		.out_empty         (),                                                                                                 // (terminated)
		.in_error          (1'b0),                                                                                             // (terminated)
		.out_error         (),                                                                                                 // (terminated)
		.in_channel        (1'b0),                                                                                             // (terminated)
		.out_channel       ()                                                                                                  // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (74),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (54),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (55),
		.PKT_TRANS_POSTED          (56),
		.PKT_TRANS_WRITE           (57),
		.PKT_TRANS_READ            (58),
		.PKT_TRANS_LOCK            (59),
		.PKT_SRC_ID_H              (79),
		.PKT_SRC_ID_L              (76),
		.PKT_DEST_ID_H             (83),
		.PKT_DEST_ID_L             (80),
		.PKT_BURSTWRAP_H           (66),
		.PKT_BURSTWRAP_L           (64),
		.PKT_BYTE_CNT_H            (63),
		.PKT_BYTE_CNT_L            (61),
		.PKT_PROTECTION_H          (87),
		.PKT_PROTECTION_L          (85),
		.PKT_RESPONSE_STATUS_H     (93),
		.PKT_RESPONSE_STATUS_L     (92),
		.PKT_BURST_SIZE_H          (69),
		.PKT_BURST_SIZE_L          (67),
		.ST_CHANNEL_W              (12),
		.ST_DATA_W                 (94),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) data_h_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                        //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                 //       clk_reset.reset
		.m0_address              (data_h_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (data_h_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (data_h_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (data_h_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (data_h_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (data_h_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (data_h_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (data_h_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (data_h_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (data_h_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (data_h_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (data_h_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (data_h_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (data_h_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (data_h_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (data_h_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src5_ready),                                                  //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src5_valid),                                                  //                .valid
		.cp_data                 (cmd_xbar_demux_001_src5_data),                                                   //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src5_startofpacket),                                          //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src5_endofpacket),                                            //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src5_channel),                                                //                .channel
		.rf_sink_ready           (data_h_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (data_h_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (data_h_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (data_h_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (data_h_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (data_h_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (data_h_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (data_h_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (data_h_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (data_h_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (data_h_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (data_h_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (data_h_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (data_h_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (data_h_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (data_h_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (95),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) data_h_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                        //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                 // clk_reset.reset
		.in_data           (data_h_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (data_h_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (data_h_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (data_h_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (data_h_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (data_h_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (data_h_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (data_h_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (data_h_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (data_h_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                          // (terminated)
		.csr_read          (1'b0),                                                                           // (terminated)
		.csr_write         (1'b0),                                                                           // (terminated)
		.csr_readdata      (),                                                                               // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                           // (terminated)
		.almost_full_data  (),                                                                               // (terminated)
		.almost_empty_data (),                                                                               // (terminated)
		.in_empty          (1'b0),                                                                           // (terminated)
		.out_empty         (),                                                                               // (terminated)
		.in_error          (1'b0),                                                                           // (terminated)
		.out_error         (),                                                                               // (terminated)
		.in_channel        (1'b0),                                                                           // (terminated)
		.out_channel       ()                                                                                // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (74),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (54),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (55),
		.PKT_TRANS_POSTED          (56),
		.PKT_TRANS_WRITE           (57),
		.PKT_TRANS_READ            (58),
		.PKT_TRANS_LOCK            (59),
		.PKT_SRC_ID_H              (79),
		.PKT_SRC_ID_L              (76),
		.PKT_DEST_ID_H             (83),
		.PKT_DEST_ID_L             (80),
		.PKT_BURSTWRAP_H           (66),
		.PKT_BURSTWRAP_L           (64),
		.PKT_BYTE_CNT_H            (63),
		.PKT_BYTE_CNT_L            (61),
		.PKT_PROTECTION_H          (87),
		.PKT_PROTECTION_L          (85),
		.PKT_RESPONSE_STATUS_H     (93),
		.PKT_RESPONSE_STATUS_L     (92),
		.PKT_BURST_SIZE_H          (69),
		.PKT_BURST_SIZE_L          (67),
		.ST_CHANNEL_W              (12),
		.ST_DATA_W                 (94),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) sysid_control_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                  //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                           //       clk_reset.reset
		.m0_address              (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src6_ready),                                                            //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src6_valid),                                                            //                .valid
		.cp_data                 (cmd_xbar_demux_001_src6_data),                                                             //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src6_startofpacket),                                                    //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src6_endofpacket),                                                      //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src6_channel),                                                          //                .channel
		.rf_sink_ready           (sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (95),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                  //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                           // clk_reset.reset
		.in_data           (sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                    // (terminated)
		.csr_read          (1'b0),                                                                                     // (terminated)
		.csr_write         (1'b0),                                                                                     // (terminated)
		.csr_readdata      (),                                                                                         // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                     // (terminated)
		.almost_full_data  (),                                                                                         // (terminated)
		.almost_empty_data (),                                                                                         // (terminated)
		.in_empty          (1'b0),                                                                                     // (terminated)
		.out_empty         (),                                                                                         // (terminated)
		.in_error          (1'b0),                                                                                     // (terminated)
		.out_error         (),                                                                                         // (terminated)
		.in_channel        (1'b0),                                                                                     // (terminated)
		.out_channel       ()                                                                                          // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (74),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (54),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (55),
		.PKT_TRANS_POSTED          (56),
		.PKT_TRANS_WRITE           (57),
		.PKT_TRANS_READ            (58),
		.PKT_TRANS_LOCK            (59),
		.PKT_SRC_ID_H              (79),
		.PKT_SRC_ID_L              (76),
		.PKT_DEST_ID_H             (83),
		.PKT_DEST_ID_L             (80),
		.PKT_BURSTWRAP_H           (66),
		.PKT_BURSTWRAP_L           (64),
		.PKT_BYTE_CNT_H            (63),
		.PKT_BYTE_CNT_L            (61),
		.PKT_PROTECTION_H          (87),
		.PKT_PROTECTION_L          (85),
		.PKT_RESPONSE_STATUS_H     (93),
		.PKT_RESPONSE_STATUS_L     (92),
		.PKT_BURST_SIZE_H          (69),
		.PKT_BURST_SIZE_L          (67),
		.ST_CHANNEL_W              (12),
		.ST_DATA_W                 (94),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) data_l_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                        //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                 //       clk_reset.reset
		.m0_address              (data_l_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (data_l_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (data_l_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (data_l_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (data_l_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (data_l_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (data_l_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (data_l_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (data_l_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (data_l_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (data_l_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (data_l_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (data_l_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (data_l_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (data_l_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (data_l_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src7_ready),                                                  //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src7_valid),                                                  //                .valid
		.cp_data                 (cmd_xbar_demux_001_src7_data),                                                   //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src7_startofpacket),                                          //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src7_endofpacket),                                            //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src7_channel),                                                //                .channel
		.rf_sink_ready           (data_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (data_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (data_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (data_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (data_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (data_l_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (data_l_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (data_l_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (data_l_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (data_l_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (data_l_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (data_l_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (data_l_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (data_l_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (data_l_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (data_l_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (95),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) data_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                        //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                 // clk_reset.reset
		.in_data           (data_l_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (data_l_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (data_l_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (data_l_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (data_l_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (data_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (data_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (data_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (data_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (data_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                          // (terminated)
		.csr_read          (1'b0),                                                                           // (terminated)
		.csr_write         (1'b0),                                                                           // (terminated)
		.csr_readdata      (),                                                                               // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                           // (terminated)
		.almost_full_data  (),                                                                               // (terminated)
		.almost_empty_data (),                                                                               // (terminated)
		.in_empty          (1'b0),                                                                           // (terminated)
		.out_empty         (),                                                                               // (terminated)
		.in_error          (1'b0),                                                                           // (terminated)
		.out_error         (),                                                                               // (terminated)
		.in_channel        (1'b0),                                                                           // (terminated)
		.out_channel       ()                                                                                // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (74),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (54),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (55),
		.PKT_TRANS_POSTED          (56),
		.PKT_TRANS_WRITE           (57),
		.PKT_TRANS_READ            (58),
		.PKT_TRANS_LOCK            (59),
		.PKT_SRC_ID_H              (79),
		.PKT_SRC_ID_L              (76),
		.PKT_DEST_ID_H             (83),
		.PKT_DEST_ID_L             (80),
		.PKT_BURSTWRAP_H           (66),
		.PKT_BURSTWRAP_L           (64),
		.PKT_BYTE_CNT_H            (63),
		.PKT_BYTE_CNT_L            (61),
		.PKT_PROTECTION_H          (87),
		.PKT_PROTECTION_L          (85),
		.PKT_RESPONSE_STATUS_H     (93),
		.PKT_RESPONSE_STATUS_L     (92),
		.PKT_BURST_SIZE_H          (69),
		.PKT_BURST_SIZE_L          (67),
		.ST_CHANNEL_W              (12),
		.ST_DATA_W                 (94),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) pre_come_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                          //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                   //       clk_reset.reset
		.m0_address              (pre_come_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (pre_come_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (pre_come_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (pre_come_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (pre_come_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (pre_come_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (pre_come_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (pre_come_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (pre_come_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (pre_come_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (pre_come_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (pre_come_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (pre_come_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (pre_come_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (pre_come_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (pre_come_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src8_ready),                                                    //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src8_valid),                                                    //                .valid
		.cp_data                 (cmd_xbar_demux_001_src8_data),                                                     //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src8_startofpacket),                                            //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src8_endofpacket),                                              //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src8_channel),                                                  //                .channel
		.rf_sink_ready           (pre_come_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (pre_come_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (pre_come_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (pre_come_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (pre_come_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (pre_come_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (pre_come_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (pre_come_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (pre_come_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (pre_come_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (pre_come_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (pre_come_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (pre_come_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (pre_come_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (pre_come_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (pre_come_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (95),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) pre_come_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                          //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                   // clk_reset.reset
		.in_data           (pre_come_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (pre_come_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (pre_come_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (pre_come_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (pre_come_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (pre_come_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (pre_come_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (pre_come_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (pre_come_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (pre_come_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                            // (terminated)
		.csr_read          (1'b0),                                                                             // (terminated)
		.csr_write         (1'b0),                                                                             // (terminated)
		.csr_readdata      (),                                                                                 // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                             // (terminated)
		.almost_full_data  (),                                                                                 // (terminated)
		.almost_empty_data (),                                                                                 // (terminated)
		.in_empty          (1'b0),                                                                             // (terminated)
		.out_empty         (),                                                                                 // (terminated)
		.in_error          (1'b0),                                                                             // (terminated)
		.out_error         (),                                                                                 // (terminated)
		.in_channel        (1'b0),                                                                             // (terminated)
		.out_channel       ()                                                                                  // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (74),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (54),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (55),
		.PKT_TRANS_POSTED          (56),
		.PKT_TRANS_WRITE           (57),
		.PKT_TRANS_READ            (58),
		.PKT_TRANS_LOCK            (59),
		.PKT_SRC_ID_H              (79),
		.PKT_SRC_ID_L              (76),
		.PKT_DEST_ID_H             (83),
		.PKT_DEST_ID_L             (80),
		.PKT_BURSTWRAP_H           (66),
		.PKT_BURSTWRAP_L           (64),
		.PKT_BYTE_CNT_H            (63),
		.PKT_BYTE_CNT_L            (61),
		.PKT_PROTECTION_H          (87),
		.PKT_PROTECTION_L          (85),
		.PKT_RESPONSE_STATUS_H     (93),
		.PKT_RESPONSE_STATUS_L     (92),
		.PKT_BURST_SIZE_H          (69),
		.PKT_BURST_SIZE_L          (67),
		.ST_CHANNEL_W              (12),
		.ST_DATA_W                 (94),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) tx_data_l_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                           //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                    //       clk_reset.reset
		.m0_address              (tx_data_l_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (tx_data_l_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (tx_data_l_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (tx_data_l_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (tx_data_l_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (tx_data_l_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (tx_data_l_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (tx_data_l_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (tx_data_l_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (tx_data_l_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (tx_data_l_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (tx_data_l_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (tx_data_l_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (tx_data_l_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (tx_data_l_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (tx_data_l_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src9_ready),                                                     //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src9_valid),                                                     //                .valid
		.cp_data                 (cmd_xbar_demux_001_src9_data),                                                      //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src9_startofpacket),                                             //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src9_endofpacket),                                               //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src9_channel),                                                   //                .channel
		.rf_sink_ready           (tx_data_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (tx_data_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (tx_data_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (tx_data_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (tx_data_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (tx_data_l_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (tx_data_l_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (tx_data_l_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (tx_data_l_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (tx_data_l_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (tx_data_l_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (tx_data_l_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (tx_data_l_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (tx_data_l_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (tx_data_l_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (tx_data_l_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (95),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) tx_data_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                           //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                    // clk_reset.reset
		.in_data           (tx_data_l_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (tx_data_l_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (tx_data_l_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (tx_data_l_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (tx_data_l_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (tx_data_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (tx_data_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (tx_data_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (tx_data_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (tx_data_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                             // (terminated)
		.csr_read          (1'b0),                                                                              // (terminated)
		.csr_write         (1'b0),                                                                              // (terminated)
		.csr_readdata      (),                                                                                  // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                              // (terminated)
		.almost_full_data  (),                                                                                  // (terminated)
		.almost_empty_data (),                                                                                  // (terminated)
		.in_empty          (1'b0),                                                                              // (terminated)
		.out_empty         (),                                                                                  // (terminated)
		.in_error          (1'b0),                                                                              // (terminated)
		.out_error         (),                                                                                  // (terminated)
		.in_channel        (1'b0),                                                                              // (terminated)
		.out_channel       ()                                                                                   // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (74),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (54),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (55),
		.PKT_TRANS_POSTED          (56),
		.PKT_TRANS_WRITE           (57),
		.PKT_TRANS_READ            (58),
		.PKT_TRANS_LOCK            (59),
		.PKT_SRC_ID_H              (79),
		.PKT_SRC_ID_L              (76),
		.PKT_DEST_ID_H             (83),
		.PKT_DEST_ID_L             (80),
		.PKT_BURSTWRAP_H           (66),
		.PKT_BURSTWRAP_L           (64),
		.PKT_BYTE_CNT_H            (63),
		.PKT_BYTE_CNT_L            (61),
		.PKT_PROTECTION_H          (87),
		.PKT_PROTECTION_L          (85),
		.PKT_RESPONSE_STATUS_H     (93),
		.PKT_RESPONSE_STATUS_L     (92),
		.PKT_BURST_SIZE_H          (69),
		.PKT_BURST_SIZE_L          (67),
		.ST_CHANNEL_W              (12),
		.ST_DATA_W                 (94),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) tx_data_h_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                           //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                    //       clk_reset.reset
		.m0_address              (tx_data_h_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (tx_data_h_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (tx_data_h_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (tx_data_h_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (tx_data_h_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (tx_data_h_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (tx_data_h_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (tx_data_h_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (tx_data_h_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (tx_data_h_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (tx_data_h_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (tx_data_h_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (tx_data_h_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (tx_data_h_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (tx_data_h_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (tx_data_h_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src10_ready),                                                    //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src10_valid),                                                    //                .valid
		.cp_data                 (cmd_xbar_demux_001_src10_data),                                                     //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src10_startofpacket),                                            //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src10_endofpacket),                                              //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src10_channel),                                                  //                .channel
		.rf_sink_ready           (tx_data_h_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (tx_data_h_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (tx_data_h_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (tx_data_h_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (tx_data_h_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (tx_data_h_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (tx_data_h_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (tx_data_h_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (tx_data_h_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (tx_data_h_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (tx_data_h_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (tx_data_h_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (tx_data_h_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (tx_data_h_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (tx_data_h_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (tx_data_h_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (95),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) tx_data_h_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                           //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                    // clk_reset.reset
		.in_data           (tx_data_h_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (tx_data_h_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (tx_data_h_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (tx_data_h_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (tx_data_h_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (tx_data_h_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (tx_data_h_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (tx_data_h_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (tx_data_h_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (tx_data_h_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                             // (terminated)
		.csr_read          (1'b0),                                                                              // (terminated)
		.csr_write         (1'b0),                                                                              // (terminated)
		.csr_readdata      (),                                                                                  // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                              // (terminated)
		.almost_full_data  (),                                                                                  // (terminated)
		.almost_empty_data (),                                                                                  // (terminated)
		.in_empty          (1'b0),                                                                              // (terminated)
		.out_empty         (),                                                                                  // (terminated)
		.in_error          (1'b0),                                                                              // (terminated)
		.out_error         (),                                                                                  // (terminated)
		.in_channel        (1'b0),                                                                              // (terminated)
		.out_channel       ()                                                                                   // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (74),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (54),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (55),
		.PKT_TRANS_POSTED          (56),
		.PKT_TRANS_WRITE           (57),
		.PKT_TRANS_READ            (58),
		.PKT_TRANS_LOCK            (59),
		.PKT_SRC_ID_H              (79),
		.PKT_SRC_ID_L              (76),
		.PKT_DEST_ID_H             (83),
		.PKT_DEST_ID_L             (80),
		.PKT_BURSTWRAP_H           (66),
		.PKT_BURSTWRAP_L           (64),
		.PKT_BYTE_CNT_H            (63),
		.PKT_BYTE_CNT_L            (61),
		.PKT_PROTECTION_H          (87),
		.PKT_PROTECTION_L          (85),
		.PKT_RESPONSE_STATUS_H     (93),
		.PKT_RESPONSE_STATUS_L     (92),
		.PKT_BURST_SIZE_H          (69),
		.PKT_BURST_SIZE_L          (67),
		.ST_CHANNEL_W              (12),
		.ST_DATA_W                 (94),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) tx_data_valid_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                               //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                        //       clk_reset.reset
		.m0_address              (tx_data_valid_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (tx_data_valid_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (tx_data_valid_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (tx_data_valid_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (tx_data_valid_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (tx_data_valid_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (tx_data_valid_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (tx_data_valid_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (tx_data_valid_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (tx_data_valid_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (tx_data_valid_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (tx_data_valid_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (tx_data_valid_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (tx_data_valid_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (tx_data_valid_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (tx_data_valid_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src11_ready),                                                        //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src11_valid),                                                        //                .valid
		.cp_data                 (cmd_xbar_demux_001_src11_data),                                                         //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src11_startofpacket),                                                //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src11_endofpacket),                                                  //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src11_channel),                                                      //                .channel
		.rf_sink_ready           (tx_data_valid_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (tx_data_valid_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (tx_data_valid_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (tx_data_valid_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (tx_data_valid_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (tx_data_valid_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (tx_data_valid_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (tx_data_valid_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (tx_data_valid_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (tx_data_valid_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (tx_data_valid_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (tx_data_valid_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (tx_data_valid_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (tx_data_valid_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (tx_data_valid_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (tx_data_valid_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (95),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) tx_data_valid_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                               //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                        // clk_reset.reset
		.in_data           (tx_data_valid_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (tx_data_valid_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (tx_data_valid_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (tx_data_valid_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (tx_data_valid_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (tx_data_valid_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (tx_data_valid_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (tx_data_valid_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (tx_data_valid_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (tx_data_valid_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                 // (terminated)
		.csr_read          (1'b0),                                                                                  // (terminated)
		.csr_write         (1'b0),                                                                                  // (terminated)
		.csr_readdata      (),                                                                                      // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                  // (terminated)
		.almost_full_data  (),                                                                                      // (terminated)
		.almost_empty_data (),                                                                                      // (terminated)
		.in_empty          (1'b0),                                                                                  // (terminated)
		.out_empty         (),                                                                                      // (terminated)
		.in_error          (1'b0),                                                                                  // (terminated)
		.out_error         (),                                                                                      // (terminated)
		.in_channel        (1'b0),                                                                                  // (terminated)
		.out_channel       ()                                                                                       // (terminated)
	);

	NIOS2_addr_router addr_router (
		.sink_ready         (cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                            //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                     // clk_reset.reset
		.src_ready          (addr_router_src_ready),                                                              //       src.ready
		.src_valid          (addr_router_src_valid),                                                              //          .valid
		.src_data           (addr_router_src_data),                                                               //          .data
		.src_channel        (addr_router_src_channel),                                                            //          .channel
		.src_startofpacket  (addr_router_src_startofpacket),                                                      //          .startofpacket
		.src_endofpacket    (addr_router_src_endofpacket)                                                         //          .endofpacket
	);

	NIOS2_addr_router_001 addr_router_001 (
		.sink_ready         (cpu_data_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (cpu_data_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (cpu_data_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (cpu_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (cpu_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                     //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                              // clk_reset.reset
		.src_ready          (addr_router_001_src_ready),                                                   //       src.ready
		.src_valid          (addr_router_001_src_valid),                                                   //          .valid
		.src_data           (addr_router_001_src_data),                                                    //          .data
		.src_channel        (addr_router_001_src_channel),                                                 //          .channel
		.src_startofpacket  (addr_router_001_src_startofpacket),                                           //          .startofpacket
		.src_endofpacket    (addr_router_001_src_endofpacket)                                              //          .endofpacket
	);

	NIOS2_id_router id_router (
		.sink_ready         (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                          //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                   // clk_reset.reset
		.src_ready          (id_router_src_ready),                                                              //       src.ready
		.src_valid          (id_router_src_valid),                                                              //          .valid
		.src_data           (id_router_src_data),                                                               //          .data
		.src_channel        (id_router_src_channel),                                                            //          .channel
		.src_startofpacket  (id_router_src_startofpacket),                                                      //          .startofpacket
		.src_endofpacket    (id_router_src_endofpacket)                                                         //          .endofpacket
	);

	NIOS2_id_router id_router_001 (
		.sink_ready         (ram_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (ram_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (ram_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (ram_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (ram_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                           //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                    // clk_reset.reset
		.src_ready          (id_router_001_src_ready),                                           //       src.ready
		.src_valid          (id_router_001_src_valid),                                           //          .valid
		.src_data           (id_router_001_src_data),                                            //          .data
		.src_channel        (id_router_001_src_channel),                                         //          .channel
		.src_startofpacket  (id_router_001_src_startofpacket),                                   //          .startofpacket
		.src_endofpacket    (id_router_001_src_endofpacket)                                      //          .endofpacket
	);

	NIOS2_id_router id_router_002 (
		.sink_ready         (epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (epcs_flash_controller_0_epcs_control_port_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                                              //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                                       // clk_reset.reset
		.src_ready          (id_router_002_src_ready),                                                                              //       src.ready
		.src_valid          (id_router_002_src_valid),                                                                              //          .valid
		.src_data           (id_router_002_src_data),                                                                               //          .data
		.src_channel        (id_router_002_src_channel),                                                                            //          .channel
		.src_startofpacket  (id_router_002_src_startofpacket),                                                                      //          .startofpacket
		.src_endofpacket    (id_router_002_src_endofpacket)                                                                         //          .endofpacket
	);

	NIOS2_id_router_003 id_router_003 (
		.sink_ready         (uart_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (uart_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (uart_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (uart_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (uart_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                            //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                     // clk_reset.reset
		.src_ready          (id_router_003_src_ready),                                            //       src.ready
		.src_valid          (id_router_003_src_valid),                                            //          .valid
		.src_data           (id_router_003_src_data),                                             //          .data
		.src_channel        (id_router_003_src_channel),                                          //          .channel
		.src_startofpacket  (id_router_003_src_startofpacket),                                    //          .startofpacket
		.src_endofpacket    (id_router_003_src_endofpacket)                                       //          .endofpacket
	);

	NIOS2_id_router_003 id_router_004 (
		.sink_ready         (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                                //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                         // clk_reset.reset
		.src_ready          (id_router_004_src_ready),                                                                //       src.ready
		.src_valid          (id_router_004_src_valid),                                                                //          .valid
		.src_data           (id_router_004_src_data),                                                                 //          .data
		.src_channel        (id_router_004_src_channel),                                                              //          .channel
		.src_startofpacket  (id_router_004_src_startofpacket),                                                        //          .startofpacket
		.src_endofpacket    (id_router_004_src_endofpacket)                                                           //          .endofpacket
	);

	NIOS2_id_router_003 id_router_005 (
		.sink_ready         (data_h_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (data_h_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (data_h_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (data_h_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (data_h_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                              //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                       // clk_reset.reset
		.src_ready          (id_router_005_src_ready),                                              //       src.ready
		.src_valid          (id_router_005_src_valid),                                              //          .valid
		.src_data           (id_router_005_src_data),                                               //          .data
		.src_channel        (id_router_005_src_channel),                                            //          .channel
		.src_startofpacket  (id_router_005_src_startofpacket),                                      //          .startofpacket
		.src_endofpacket    (id_router_005_src_endofpacket)                                         //          .endofpacket
	);

	NIOS2_id_router_003 id_router_006 (
		.sink_ready         (sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                        //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                 // clk_reset.reset
		.src_ready          (id_router_006_src_ready),                                                        //       src.ready
		.src_valid          (id_router_006_src_valid),                                                        //          .valid
		.src_data           (id_router_006_src_data),                                                         //          .data
		.src_channel        (id_router_006_src_channel),                                                      //          .channel
		.src_startofpacket  (id_router_006_src_startofpacket),                                                //          .startofpacket
		.src_endofpacket    (id_router_006_src_endofpacket)                                                   //          .endofpacket
	);

	NIOS2_id_router_003 id_router_007 (
		.sink_ready         (data_l_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (data_l_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (data_l_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (data_l_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (data_l_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                              //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                       // clk_reset.reset
		.src_ready          (id_router_007_src_ready),                                              //       src.ready
		.src_valid          (id_router_007_src_valid),                                              //          .valid
		.src_data           (id_router_007_src_data),                                               //          .data
		.src_channel        (id_router_007_src_channel),                                            //          .channel
		.src_startofpacket  (id_router_007_src_startofpacket),                                      //          .startofpacket
		.src_endofpacket    (id_router_007_src_endofpacket)                                         //          .endofpacket
	);

	NIOS2_id_router_003 id_router_008 (
		.sink_ready         (pre_come_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (pre_come_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (pre_come_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (pre_come_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (pre_come_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                         // clk_reset.reset
		.src_ready          (id_router_008_src_ready),                                                //       src.ready
		.src_valid          (id_router_008_src_valid),                                                //          .valid
		.src_data           (id_router_008_src_data),                                                 //          .data
		.src_channel        (id_router_008_src_channel),                                              //          .channel
		.src_startofpacket  (id_router_008_src_startofpacket),                                        //          .startofpacket
		.src_endofpacket    (id_router_008_src_endofpacket)                                           //          .endofpacket
	);

	NIOS2_id_router_003 id_router_009 (
		.sink_ready         (tx_data_l_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (tx_data_l_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (tx_data_l_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (tx_data_l_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (tx_data_l_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                 //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                          // clk_reset.reset
		.src_ready          (id_router_009_src_ready),                                                 //       src.ready
		.src_valid          (id_router_009_src_valid),                                                 //          .valid
		.src_data           (id_router_009_src_data),                                                  //          .data
		.src_channel        (id_router_009_src_channel),                                               //          .channel
		.src_startofpacket  (id_router_009_src_startofpacket),                                         //          .startofpacket
		.src_endofpacket    (id_router_009_src_endofpacket)                                            //          .endofpacket
	);

	NIOS2_id_router_003 id_router_010 (
		.sink_ready         (tx_data_h_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (tx_data_h_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (tx_data_h_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (tx_data_h_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (tx_data_h_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                 //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                          // clk_reset.reset
		.src_ready          (id_router_010_src_ready),                                                 //       src.ready
		.src_valid          (id_router_010_src_valid),                                                 //          .valid
		.src_data           (id_router_010_src_data),                                                  //          .data
		.src_channel        (id_router_010_src_channel),                                               //          .channel
		.src_startofpacket  (id_router_010_src_startofpacket),                                         //          .startofpacket
		.src_endofpacket    (id_router_010_src_endofpacket)                                            //          .endofpacket
	);

	NIOS2_id_router_003 id_router_011 (
		.sink_ready         (tx_data_valid_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (tx_data_valid_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (tx_data_valid_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (tx_data_valid_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (tx_data_valid_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                     //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                              // clk_reset.reset
		.src_ready          (id_router_011_src_ready),                                                     //       src.ready
		.src_valid          (id_router_011_src_valid),                                                     //          .valid
		.src_data           (id_router_011_src_data),                                                      //          .data
		.src_channel        (id_router_011_src_channel),                                                   //          .channel
		.src_startofpacket  (id_router_011_src_startofpacket),                                             //          .startofpacket
		.src_endofpacket    (id_router_011_src_endofpacket)                                                //          .endofpacket
	);

	altera_merlin_traffic_limiter #(
		.PKT_DEST_ID_H             (83),
		.PKT_DEST_ID_L             (80),
		.PKT_TRANS_POSTED          (56),
		.PKT_TRANS_WRITE           (57),
		.MAX_OUTSTANDING_RESPONSES (1),
		.PIPELINED                 (0),
		.ST_DATA_W                 (94),
		.ST_CHANNEL_W              (12),
		.VALID_WIDTH               (12),
		.ENFORCE_ORDER             (1),
		.PREVENT_HAZARDS           (0),
		.PKT_BYTE_CNT_H            (63),
		.PKT_BYTE_CNT_L            (61),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32)
	) limiter (
		.clk                    (clk_clk),                        //       clk.clk
		.reset                  (rst_controller_reset_out_reset), // clk_reset.reset
		.cmd_sink_ready         (addr_router_src_ready),          //  cmd_sink.ready
		.cmd_sink_valid         (addr_router_src_valid),          //          .valid
		.cmd_sink_data          (addr_router_src_data),           //          .data
		.cmd_sink_channel       (addr_router_src_channel),        //          .channel
		.cmd_sink_startofpacket (addr_router_src_startofpacket),  //          .startofpacket
		.cmd_sink_endofpacket   (addr_router_src_endofpacket),    //          .endofpacket
		.cmd_src_ready          (limiter_cmd_src_ready),          //   cmd_src.ready
		.cmd_src_data           (limiter_cmd_src_data),           //          .data
		.cmd_src_channel        (limiter_cmd_src_channel),        //          .channel
		.cmd_src_startofpacket  (limiter_cmd_src_startofpacket),  //          .startofpacket
		.cmd_src_endofpacket    (limiter_cmd_src_endofpacket),    //          .endofpacket
		.rsp_sink_ready         (rsp_xbar_mux_src_ready),         //  rsp_sink.ready
		.rsp_sink_valid         (rsp_xbar_mux_src_valid),         //          .valid
		.rsp_sink_channel       (rsp_xbar_mux_src_channel),       //          .channel
		.rsp_sink_data          (rsp_xbar_mux_src_data),          //          .data
		.rsp_sink_startofpacket (rsp_xbar_mux_src_startofpacket), //          .startofpacket
		.rsp_sink_endofpacket   (rsp_xbar_mux_src_endofpacket),   //          .endofpacket
		.rsp_src_ready          (limiter_rsp_src_ready),          //   rsp_src.ready
		.rsp_src_valid          (limiter_rsp_src_valid),          //          .valid
		.rsp_src_data           (limiter_rsp_src_data),           //          .data
		.rsp_src_channel        (limiter_rsp_src_channel),        //          .channel
		.rsp_src_startofpacket  (limiter_rsp_src_startofpacket),  //          .startofpacket
		.rsp_src_endofpacket    (limiter_rsp_src_endofpacket),    //          .endofpacket
		.cmd_src_valid          (limiter_cmd_valid_data)          // cmd_valid.data
	);

	altera_merlin_traffic_limiter #(
		.PKT_DEST_ID_H             (83),
		.PKT_DEST_ID_L             (80),
		.PKT_TRANS_POSTED          (56),
		.PKT_TRANS_WRITE           (57),
		.MAX_OUTSTANDING_RESPONSES (1),
		.PIPELINED                 (0),
		.ST_DATA_W                 (94),
		.ST_CHANNEL_W              (12),
		.VALID_WIDTH               (12),
		.ENFORCE_ORDER             (1),
		.PREVENT_HAZARDS           (0),
		.PKT_BYTE_CNT_H            (63),
		.PKT_BYTE_CNT_L            (61),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32)
	) limiter_001 (
		.clk                    (clk_clk),                            //       clk.clk
		.reset                  (rst_controller_reset_out_reset),     // clk_reset.reset
		.cmd_sink_ready         (addr_router_001_src_ready),          //  cmd_sink.ready
		.cmd_sink_valid         (addr_router_001_src_valid),          //          .valid
		.cmd_sink_data          (addr_router_001_src_data),           //          .data
		.cmd_sink_channel       (addr_router_001_src_channel),        //          .channel
		.cmd_sink_startofpacket (addr_router_001_src_startofpacket),  //          .startofpacket
		.cmd_sink_endofpacket   (addr_router_001_src_endofpacket),    //          .endofpacket
		.cmd_src_ready          (limiter_001_cmd_src_ready),          //   cmd_src.ready
		.cmd_src_data           (limiter_001_cmd_src_data),           //          .data
		.cmd_src_channel        (limiter_001_cmd_src_channel),        //          .channel
		.cmd_src_startofpacket  (limiter_001_cmd_src_startofpacket),  //          .startofpacket
		.cmd_src_endofpacket    (limiter_001_cmd_src_endofpacket),    //          .endofpacket
		.rsp_sink_ready         (rsp_xbar_mux_001_src_ready),         //  rsp_sink.ready
		.rsp_sink_valid         (rsp_xbar_mux_001_src_valid),         //          .valid
		.rsp_sink_channel       (rsp_xbar_mux_001_src_channel),       //          .channel
		.rsp_sink_data          (rsp_xbar_mux_001_src_data),          //          .data
		.rsp_sink_startofpacket (rsp_xbar_mux_001_src_startofpacket), //          .startofpacket
		.rsp_sink_endofpacket   (rsp_xbar_mux_001_src_endofpacket),   //          .endofpacket
		.rsp_src_ready          (limiter_001_rsp_src_ready),          //   rsp_src.ready
		.rsp_src_valid          (limiter_001_rsp_src_valid),          //          .valid
		.rsp_src_data           (limiter_001_rsp_src_data),           //          .data
		.rsp_src_channel        (limiter_001_rsp_src_channel),        //          .channel
		.rsp_src_startofpacket  (limiter_001_rsp_src_startofpacket),  //          .startofpacket
		.rsp_src_endofpacket    (limiter_001_rsp_src_endofpacket),    //          .endofpacket
		.cmd_src_valid          (limiter_001_cmd_valid_data)          // cmd_valid.data
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (2),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2)
	) rst_controller (
		.reset_in0  (~reset_reset_n),                    // reset_in0.reset
		.reset_in1  (cpu_jtag_debug_module_reset_reset), // reset_in1.reset
		.clk        (clk_clk),                           //       clk.clk
		.reset_out  (rst_controller_reset_out_reset),    // reset_out.reset
		.reset_in2  (1'b0),                              // (terminated)
		.reset_in3  (1'b0),                              // (terminated)
		.reset_in4  (1'b0),                              // (terminated)
		.reset_in5  (1'b0),                              // (terminated)
		.reset_in6  (1'b0),                              // (terminated)
		.reset_in7  (1'b0),                              // (terminated)
		.reset_in8  (1'b0),                              // (terminated)
		.reset_in9  (1'b0),                              // (terminated)
		.reset_in10 (1'b0),                              // (terminated)
		.reset_in11 (1'b0),                              // (terminated)
		.reset_in12 (1'b0),                              // (terminated)
		.reset_in13 (1'b0),                              // (terminated)
		.reset_in14 (1'b0),                              // (terminated)
		.reset_in15 (1'b0)                               // (terminated)
	);

	NIOS2_cmd_xbar_demux cmd_xbar_demux (
		.clk                (clk_clk),                           //        clk.clk
		.reset              (rst_controller_reset_out_reset),    //  clk_reset.reset
		.sink_ready         (limiter_cmd_src_ready),             //       sink.ready
		.sink_channel       (limiter_cmd_src_channel),           //           .channel
		.sink_data          (limiter_cmd_src_data),              //           .data
		.sink_startofpacket (limiter_cmd_src_startofpacket),     //           .startofpacket
		.sink_endofpacket   (limiter_cmd_src_endofpacket),       //           .endofpacket
		.sink_valid         (limiter_cmd_valid_data),            // sink_valid.data
		.src0_ready         (cmd_xbar_demux_src0_ready),         //       src0.ready
		.src0_valid         (cmd_xbar_demux_src0_valid),         //           .valid
		.src0_data          (cmd_xbar_demux_src0_data),          //           .data
		.src0_channel       (cmd_xbar_demux_src0_channel),       //           .channel
		.src0_startofpacket (cmd_xbar_demux_src0_startofpacket), //           .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_src0_endofpacket),   //           .endofpacket
		.src1_ready         (cmd_xbar_demux_src1_ready),         //       src1.ready
		.src1_valid         (cmd_xbar_demux_src1_valid),         //           .valid
		.src1_data          (cmd_xbar_demux_src1_data),          //           .data
		.src1_channel       (cmd_xbar_demux_src1_channel),       //           .channel
		.src1_startofpacket (cmd_xbar_demux_src1_startofpacket), //           .startofpacket
		.src1_endofpacket   (cmd_xbar_demux_src1_endofpacket),   //           .endofpacket
		.src2_ready         (cmd_xbar_demux_src2_ready),         //       src2.ready
		.src2_valid         (cmd_xbar_demux_src2_valid),         //           .valid
		.src2_data          (cmd_xbar_demux_src2_data),          //           .data
		.src2_channel       (cmd_xbar_demux_src2_channel),       //           .channel
		.src2_startofpacket (cmd_xbar_demux_src2_startofpacket), //           .startofpacket
		.src2_endofpacket   (cmd_xbar_demux_src2_endofpacket)    //           .endofpacket
	);

	NIOS2_cmd_xbar_demux_001 cmd_xbar_demux_001 (
		.clk                 (clk_clk),                                //        clk.clk
		.reset               (rst_controller_reset_out_reset),         //  clk_reset.reset
		.sink_ready          (limiter_001_cmd_src_ready),              //       sink.ready
		.sink_channel        (limiter_001_cmd_src_channel),            //           .channel
		.sink_data           (limiter_001_cmd_src_data),               //           .data
		.sink_startofpacket  (limiter_001_cmd_src_startofpacket),      //           .startofpacket
		.sink_endofpacket    (limiter_001_cmd_src_endofpacket),        //           .endofpacket
		.sink_valid          (limiter_001_cmd_valid_data),             // sink_valid.data
		.src0_ready          (cmd_xbar_demux_001_src0_ready),          //       src0.ready
		.src0_valid          (cmd_xbar_demux_001_src0_valid),          //           .valid
		.src0_data           (cmd_xbar_demux_001_src0_data),           //           .data
		.src0_channel        (cmd_xbar_demux_001_src0_channel),        //           .channel
		.src0_startofpacket  (cmd_xbar_demux_001_src0_startofpacket),  //           .startofpacket
		.src0_endofpacket    (cmd_xbar_demux_001_src0_endofpacket),    //           .endofpacket
		.src1_ready          (cmd_xbar_demux_001_src1_ready),          //       src1.ready
		.src1_valid          (cmd_xbar_demux_001_src1_valid),          //           .valid
		.src1_data           (cmd_xbar_demux_001_src1_data),           //           .data
		.src1_channel        (cmd_xbar_demux_001_src1_channel),        //           .channel
		.src1_startofpacket  (cmd_xbar_demux_001_src1_startofpacket),  //           .startofpacket
		.src1_endofpacket    (cmd_xbar_demux_001_src1_endofpacket),    //           .endofpacket
		.src2_ready          (cmd_xbar_demux_001_src2_ready),          //       src2.ready
		.src2_valid          (cmd_xbar_demux_001_src2_valid),          //           .valid
		.src2_data           (cmd_xbar_demux_001_src2_data),           //           .data
		.src2_channel        (cmd_xbar_demux_001_src2_channel),        //           .channel
		.src2_startofpacket  (cmd_xbar_demux_001_src2_startofpacket),  //           .startofpacket
		.src2_endofpacket    (cmd_xbar_demux_001_src2_endofpacket),    //           .endofpacket
		.src3_ready          (cmd_xbar_demux_001_src3_ready),          //       src3.ready
		.src3_valid          (cmd_xbar_demux_001_src3_valid),          //           .valid
		.src3_data           (cmd_xbar_demux_001_src3_data),           //           .data
		.src3_channel        (cmd_xbar_demux_001_src3_channel),        //           .channel
		.src3_startofpacket  (cmd_xbar_demux_001_src3_startofpacket),  //           .startofpacket
		.src3_endofpacket    (cmd_xbar_demux_001_src3_endofpacket),    //           .endofpacket
		.src4_ready          (cmd_xbar_demux_001_src4_ready),          //       src4.ready
		.src4_valid          (cmd_xbar_demux_001_src4_valid),          //           .valid
		.src4_data           (cmd_xbar_demux_001_src4_data),           //           .data
		.src4_channel        (cmd_xbar_demux_001_src4_channel),        //           .channel
		.src4_startofpacket  (cmd_xbar_demux_001_src4_startofpacket),  //           .startofpacket
		.src4_endofpacket    (cmd_xbar_demux_001_src4_endofpacket),    //           .endofpacket
		.src5_ready          (cmd_xbar_demux_001_src5_ready),          //       src5.ready
		.src5_valid          (cmd_xbar_demux_001_src5_valid),          //           .valid
		.src5_data           (cmd_xbar_demux_001_src5_data),           //           .data
		.src5_channel        (cmd_xbar_demux_001_src5_channel),        //           .channel
		.src5_startofpacket  (cmd_xbar_demux_001_src5_startofpacket),  //           .startofpacket
		.src5_endofpacket    (cmd_xbar_demux_001_src5_endofpacket),    //           .endofpacket
		.src6_ready          (cmd_xbar_demux_001_src6_ready),          //       src6.ready
		.src6_valid          (cmd_xbar_demux_001_src6_valid),          //           .valid
		.src6_data           (cmd_xbar_demux_001_src6_data),           //           .data
		.src6_channel        (cmd_xbar_demux_001_src6_channel),        //           .channel
		.src6_startofpacket  (cmd_xbar_demux_001_src6_startofpacket),  //           .startofpacket
		.src6_endofpacket    (cmd_xbar_demux_001_src6_endofpacket),    //           .endofpacket
		.src7_ready          (cmd_xbar_demux_001_src7_ready),          //       src7.ready
		.src7_valid          (cmd_xbar_demux_001_src7_valid),          //           .valid
		.src7_data           (cmd_xbar_demux_001_src7_data),           //           .data
		.src7_channel        (cmd_xbar_demux_001_src7_channel),        //           .channel
		.src7_startofpacket  (cmd_xbar_demux_001_src7_startofpacket),  //           .startofpacket
		.src7_endofpacket    (cmd_xbar_demux_001_src7_endofpacket),    //           .endofpacket
		.src8_ready          (cmd_xbar_demux_001_src8_ready),          //       src8.ready
		.src8_valid          (cmd_xbar_demux_001_src8_valid),          //           .valid
		.src8_data           (cmd_xbar_demux_001_src8_data),           //           .data
		.src8_channel        (cmd_xbar_demux_001_src8_channel),        //           .channel
		.src8_startofpacket  (cmd_xbar_demux_001_src8_startofpacket),  //           .startofpacket
		.src8_endofpacket    (cmd_xbar_demux_001_src8_endofpacket),    //           .endofpacket
		.src9_ready          (cmd_xbar_demux_001_src9_ready),          //       src9.ready
		.src9_valid          (cmd_xbar_demux_001_src9_valid),          //           .valid
		.src9_data           (cmd_xbar_demux_001_src9_data),           //           .data
		.src9_channel        (cmd_xbar_demux_001_src9_channel),        //           .channel
		.src9_startofpacket  (cmd_xbar_demux_001_src9_startofpacket),  //           .startofpacket
		.src9_endofpacket    (cmd_xbar_demux_001_src9_endofpacket),    //           .endofpacket
		.src10_ready         (cmd_xbar_demux_001_src10_ready),         //      src10.ready
		.src10_valid         (cmd_xbar_demux_001_src10_valid),         //           .valid
		.src10_data          (cmd_xbar_demux_001_src10_data),          //           .data
		.src10_channel       (cmd_xbar_demux_001_src10_channel),       //           .channel
		.src10_startofpacket (cmd_xbar_demux_001_src10_startofpacket), //           .startofpacket
		.src10_endofpacket   (cmd_xbar_demux_001_src10_endofpacket),   //           .endofpacket
		.src11_ready         (cmd_xbar_demux_001_src11_ready),         //      src11.ready
		.src11_valid         (cmd_xbar_demux_001_src11_valid),         //           .valid
		.src11_data          (cmd_xbar_demux_001_src11_data),          //           .data
		.src11_channel       (cmd_xbar_demux_001_src11_channel),       //           .channel
		.src11_startofpacket (cmd_xbar_demux_001_src11_startofpacket), //           .startofpacket
		.src11_endofpacket   (cmd_xbar_demux_001_src11_endofpacket)    //           .endofpacket
	);

	NIOS2_cmd_xbar_mux cmd_xbar_mux (
		.clk                 (clk_clk),                               //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (cmd_xbar_mux_src_ready),                //       src.ready
		.src_valid           (cmd_xbar_mux_src_valid),                //          .valid
		.src_data            (cmd_xbar_mux_src_data),                 //          .data
		.src_channel         (cmd_xbar_mux_src_channel),              //          .channel
		.src_startofpacket   (cmd_xbar_mux_src_startofpacket),        //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_src_endofpacket),          //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src0_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src0_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src0_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src0_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src0_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src0_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src0_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src0_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src0_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src0_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src0_endofpacket)    //          .endofpacket
	);

	NIOS2_cmd_xbar_mux cmd_xbar_mux_001 (
		.clk                 (clk_clk),                               //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (cmd_xbar_mux_001_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_001_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_001_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_001_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_001_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_001_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src1_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src1_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src1_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src1_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src1_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src1_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src1_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src1_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src1_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src1_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src1_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src1_endofpacket)    //          .endofpacket
	);

	NIOS2_cmd_xbar_mux cmd_xbar_mux_002 (
		.clk                 (clk_clk),                               //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (cmd_xbar_mux_002_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_002_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_002_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_002_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_002_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_002_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src2_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src2_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src2_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src2_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src2_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src2_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src2_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src2_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src2_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src2_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src2_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src2_endofpacket)    //          .endofpacket
	);

	NIOS2_rsp_xbar_demux rsp_xbar_demux (
		.clk                (clk_clk),                           //       clk.clk
		.reset              (rst_controller_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_src_ready),               //      sink.ready
		.sink_channel       (id_router_src_channel),             //          .channel
		.sink_data          (id_router_src_data),                //          .data
		.sink_startofpacket (id_router_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_src1_endofpacket)    //          .endofpacket
	);

	NIOS2_rsp_xbar_demux rsp_xbar_demux_001 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_001_src_ready),               //      sink.ready
		.sink_channel       (id_router_001_src_channel),             //          .channel
		.sink_data          (id_router_001_src_data),                //          .data
		.sink_startofpacket (id_router_001_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_001_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_001_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_001_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_001_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_001_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_001_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_001_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_001_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_001_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_001_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_001_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_001_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_001_src1_endofpacket)    //          .endofpacket
	);

	NIOS2_rsp_xbar_demux rsp_xbar_demux_002 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_002_src_ready),               //      sink.ready
		.sink_channel       (id_router_002_src_channel),             //          .channel
		.sink_data          (id_router_002_src_data),                //          .data
		.sink_startofpacket (id_router_002_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_002_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_002_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_002_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_002_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_002_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_002_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_002_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_002_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_002_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_002_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_002_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_002_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_002_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_002_src1_endofpacket)    //          .endofpacket
	);

	NIOS2_rsp_xbar_demux_003 rsp_xbar_demux_003 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_003_src_ready),               //      sink.ready
		.sink_channel       (id_router_003_src_channel),             //          .channel
		.sink_data          (id_router_003_src_data),                //          .data
		.sink_startofpacket (id_router_003_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_003_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_003_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_003_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_003_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_003_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_003_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_003_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_003_src0_endofpacket)    //          .endofpacket
	);

	NIOS2_rsp_xbar_demux_003 rsp_xbar_demux_004 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_004_src_ready),               //      sink.ready
		.sink_channel       (id_router_004_src_channel),             //          .channel
		.sink_data          (id_router_004_src_data),                //          .data
		.sink_startofpacket (id_router_004_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_004_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_004_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_004_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_004_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_004_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_004_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_004_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_004_src0_endofpacket)    //          .endofpacket
	);

	NIOS2_rsp_xbar_demux_003 rsp_xbar_demux_005 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_005_src_ready),               //      sink.ready
		.sink_channel       (id_router_005_src_channel),             //          .channel
		.sink_data          (id_router_005_src_data),                //          .data
		.sink_startofpacket (id_router_005_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_005_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_005_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_005_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_005_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_005_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_005_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_005_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_005_src0_endofpacket)    //          .endofpacket
	);

	NIOS2_rsp_xbar_demux_003 rsp_xbar_demux_006 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_006_src_ready),               //      sink.ready
		.sink_channel       (id_router_006_src_channel),             //          .channel
		.sink_data          (id_router_006_src_data),                //          .data
		.sink_startofpacket (id_router_006_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_006_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_006_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_006_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_006_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_006_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_006_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_006_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_006_src0_endofpacket)    //          .endofpacket
	);

	NIOS2_rsp_xbar_demux_003 rsp_xbar_demux_007 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_007_src_ready),               //      sink.ready
		.sink_channel       (id_router_007_src_channel),             //          .channel
		.sink_data          (id_router_007_src_data),                //          .data
		.sink_startofpacket (id_router_007_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_007_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_007_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_007_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_007_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_007_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_007_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_007_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_007_src0_endofpacket)    //          .endofpacket
	);

	NIOS2_rsp_xbar_demux_003 rsp_xbar_demux_008 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_008_src_ready),               //      sink.ready
		.sink_channel       (id_router_008_src_channel),             //          .channel
		.sink_data          (id_router_008_src_data),                //          .data
		.sink_startofpacket (id_router_008_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_008_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_008_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_008_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_008_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_008_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_008_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_008_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_008_src0_endofpacket)    //          .endofpacket
	);

	NIOS2_rsp_xbar_demux_003 rsp_xbar_demux_009 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_009_src_ready),               //      sink.ready
		.sink_channel       (id_router_009_src_channel),             //          .channel
		.sink_data          (id_router_009_src_data),                //          .data
		.sink_startofpacket (id_router_009_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_009_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_009_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_009_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_009_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_009_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_009_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_009_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_009_src0_endofpacket)    //          .endofpacket
	);

	NIOS2_rsp_xbar_demux_003 rsp_xbar_demux_010 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_010_src_ready),               //      sink.ready
		.sink_channel       (id_router_010_src_channel),             //          .channel
		.sink_data          (id_router_010_src_data),                //          .data
		.sink_startofpacket (id_router_010_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_010_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_010_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_010_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_010_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_010_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_010_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_010_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_010_src0_endofpacket)    //          .endofpacket
	);

	NIOS2_rsp_xbar_demux_003 rsp_xbar_demux_011 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_011_src_ready),               //      sink.ready
		.sink_channel       (id_router_011_src_channel),             //          .channel
		.sink_data          (id_router_011_src_data),                //          .data
		.sink_startofpacket (id_router_011_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_011_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_011_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_011_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_011_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_011_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_011_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_011_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_011_src0_endofpacket)    //          .endofpacket
	);

	NIOS2_rsp_xbar_mux rsp_xbar_mux (
		.clk                 (clk_clk),                               //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (rsp_xbar_mux_src_ready),                //       src.ready
		.src_valid           (rsp_xbar_mux_src_valid),                //          .valid
		.src_data            (rsp_xbar_mux_src_data),                 //          .data
		.src_channel         (rsp_xbar_mux_src_channel),              //          .channel
		.src_startofpacket   (rsp_xbar_mux_src_startofpacket),        //          .startofpacket
		.src_endofpacket     (rsp_xbar_mux_src_endofpacket),          //          .endofpacket
		.sink0_ready         (rsp_xbar_demux_src0_ready),             //     sink0.ready
		.sink0_valid         (rsp_xbar_demux_src0_valid),             //          .valid
		.sink0_channel       (rsp_xbar_demux_src0_channel),           //          .channel
		.sink0_data          (rsp_xbar_demux_src0_data),              //          .data
		.sink0_startofpacket (rsp_xbar_demux_src0_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (rsp_xbar_demux_src0_endofpacket),       //          .endofpacket
		.sink1_ready         (rsp_xbar_demux_001_src0_ready),         //     sink1.ready
		.sink1_valid         (rsp_xbar_demux_001_src0_valid),         //          .valid
		.sink1_channel       (rsp_xbar_demux_001_src0_channel),       //          .channel
		.sink1_data          (rsp_xbar_demux_001_src0_data),          //          .data
		.sink1_startofpacket (rsp_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.sink1_endofpacket   (rsp_xbar_demux_001_src0_endofpacket),   //          .endofpacket
		.sink2_ready         (rsp_xbar_demux_002_src0_ready),         //     sink2.ready
		.sink2_valid         (rsp_xbar_demux_002_src0_valid),         //          .valid
		.sink2_channel       (rsp_xbar_demux_002_src0_channel),       //          .channel
		.sink2_data          (rsp_xbar_demux_002_src0_data),          //          .data
		.sink2_startofpacket (rsp_xbar_demux_002_src0_startofpacket), //          .startofpacket
		.sink2_endofpacket   (rsp_xbar_demux_002_src0_endofpacket)    //          .endofpacket
	);

	NIOS2_rsp_xbar_mux_001 rsp_xbar_mux_001 (
		.clk                  (clk_clk),                               //       clk.clk
		.reset                (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready            (rsp_xbar_mux_001_src_ready),            //       src.ready
		.src_valid            (rsp_xbar_mux_001_src_valid),            //          .valid
		.src_data             (rsp_xbar_mux_001_src_data),             //          .data
		.src_channel          (rsp_xbar_mux_001_src_channel),          //          .channel
		.src_startofpacket    (rsp_xbar_mux_001_src_startofpacket),    //          .startofpacket
		.src_endofpacket      (rsp_xbar_mux_001_src_endofpacket),      //          .endofpacket
		.sink0_ready          (rsp_xbar_demux_src1_ready),             //     sink0.ready
		.sink0_valid          (rsp_xbar_demux_src1_valid),             //          .valid
		.sink0_channel        (rsp_xbar_demux_src1_channel),           //          .channel
		.sink0_data           (rsp_xbar_demux_src1_data),              //          .data
		.sink0_startofpacket  (rsp_xbar_demux_src1_startofpacket),     //          .startofpacket
		.sink0_endofpacket    (rsp_xbar_demux_src1_endofpacket),       //          .endofpacket
		.sink1_ready          (rsp_xbar_demux_001_src1_ready),         //     sink1.ready
		.sink1_valid          (rsp_xbar_demux_001_src1_valid),         //          .valid
		.sink1_channel        (rsp_xbar_demux_001_src1_channel),       //          .channel
		.sink1_data           (rsp_xbar_demux_001_src1_data),          //          .data
		.sink1_startofpacket  (rsp_xbar_demux_001_src1_startofpacket), //          .startofpacket
		.sink1_endofpacket    (rsp_xbar_demux_001_src1_endofpacket),   //          .endofpacket
		.sink2_ready          (rsp_xbar_demux_002_src1_ready),         //     sink2.ready
		.sink2_valid          (rsp_xbar_demux_002_src1_valid),         //          .valid
		.sink2_channel        (rsp_xbar_demux_002_src1_channel),       //          .channel
		.sink2_data           (rsp_xbar_demux_002_src1_data),          //          .data
		.sink2_startofpacket  (rsp_xbar_demux_002_src1_startofpacket), //          .startofpacket
		.sink2_endofpacket    (rsp_xbar_demux_002_src1_endofpacket),   //          .endofpacket
		.sink3_ready          (rsp_xbar_demux_003_src0_ready),         //     sink3.ready
		.sink3_valid          (rsp_xbar_demux_003_src0_valid),         //          .valid
		.sink3_channel        (rsp_xbar_demux_003_src0_channel),       //          .channel
		.sink3_data           (rsp_xbar_demux_003_src0_data),          //          .data
		.sink3_startofpacket  (rsp_xbar_demux_003_src0_startofpacket), //          .startofpacket
		.sink3_endofpacket    (rsp_xbar_demux_003_src0_endofpacket),   //          .endofpacket
		.sink4_ready          (rsp_xbar_demux_004_src0_ready),         //     sink4.ready
		.sink4_valid          (rsp_xbar_demux_004_src0_valid),         //          .valid
		.sink4_channel        (rsp_xbar_demux_004_src0_channel),       //          .channel
		.sink4_data           (rsp_xbar_demux_004_src0_data),          //          .data
		.sink4_startofpacket  (rsp_xbar_demux_004_src0_startofpacket), //          .startofpacket
		.sink4_endofpacket    (rsp_xbar_demux_004_src0_endofpacket),   //          .endofpacket
		.sink5_ready          (rsp_xbar_demux_005_src0_ready),         //     sink5.ready
		.sink5_valid          (rsp_xbar_demux_005_src0_valid),         //          .valid
		.sink5_channel        (rsp_xbar_demux_005_src0_channel),       //          .channel
		.sink5_data           (rsp_xbar_demux_005_src0_data),          //          .data
		.sink5_startofpacket  (rsp_xbar_demux_005_src0_startofpacket), //          .startofpacket
		.sink5_endofpacket    (rsp_xbar_demux_005_src0_endofpacket),   //          .endofpacket
		.sink6_ready          (rsp_xbar_demux_006_src0_ready),         //     sink6.ready
		.sink6_valid          (rsp_xbar_demux_006_src0_valid),         //          .valid
		.sink6_channel        (rsp_xbar_demux_006_src0_channel),       //          .channel
		.sink6_data           (rsp_xbar_demux_006_src0_data),          //          .data
		.sink6_startofpacket  (rsp_xbar_demux_006_src0_startofpacket), //          .startofpacket
		.sink6_endofpacket    (rsp_xbar_demux_006_src0_endofpacket),   //          .endofpacket
		.sink7_ready          (rsp_xbar_demux_007_src0_ready),         //     sink7.ready
		.sink7_valid          (rsp_xbar_demux_007_src0_valid),         //          .valid
		.sink7_channel        (rsp_xbar_demux_007_src0_channel),       //          .channel
		.sink7_data           (rsp_xbar_demux_007_src0_data),          //          .data
		.sink7_startofpacket  (rsp_xbar_demux_007_src0_startofpacket), //          .startofpacket
		.sink7_endofpacket    (rsp_xbar_demux_007_src0_endofpacket),   //          .endofpacket
		.sink8_ready          (rsp_xbar_demux_008_src0_ready),         //     sink8.ready
		.sink8_valid          (rsp_xbar_demux_008_src0_valid),         //          .valid
		.sink8_channel        (rsp_xbar_demux_008_src0_channel),       //          .channel
		.sink8_data           (rsp_xbar_demux_008_src0_data),          //          .data
		.sink8_startofpacket  (rsp_xbar_demux_008_src0_startofpacket), //          .startofpacket
		.sink8_endofpacket    (rsp_xbar_demux_008_src0_endofpacket),   //          .endofpacket
		.sink9_ready          (rsp_xbar_demux_009_src0_ready),         //     sink9.ready
		.sink9_valid          (rsp_xbar_demux_009_src0_valid),         //          .valid
		.sink9_channel        (rsp_xbar_demux_009_src0_channel),       //          .channel
		.sink9_data           (rsp_xbar_demux_009_src0_data),          //          .data
		.sink9_startofpacket  (rsp_xbar_demux_009_src0_startofpacket), //          .startofpacket
		.sink9_endofpacket    (rsp_xbar_demux_009_src0_endofpacket),   //          .endofpacket
		.sink10_ready         (rsp_xbar_demux_010_src0_ready),         //    sink10.ready
		.sink10_valid         (rsp_xbar_demux_010_src0_valid),         //          .valid
		.sink10_channel       (rsp_xbar_demux_010_src0_channel),       //          .channel
		.sink10_data          (rsp_xbar_demux_010_src0_data),          //          .data
		.sink10_startofpacket (rsp_xbar_demux_010_src0_startofpacket), //          .startofpacket
		.sink10_endofpacket   (rsp_xbar_demux_010_src0_endofpacket),   //          .endofpacket
		.sink11_ready         (rsp_xbar_demux_011_src0_ready),         //    sink11.ready
		.sink11_valid         (rsp_xbar_demux_011_src0_valid),         //          .valid
		.sink11_channel       (rsp_xbar_demux_011_src0_channel),       //          .channel
		.sink11_data          (rsp_xbar_demux_011_src0_data),          //          .data
		.sink11_startofpacket (rsp_xbar_demux_011_src0_startofpacket), //          .startofpacket
		.sink11_endofpacket   (rsp_xbar_demux_011_src0_endofpacket)    //          .endofpacket
	);

	NIOS2_irq_mapper irq_mapper (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),       // receiver2.irq
		.receiver3_irq (irq_mapper_receiver3_irq),       // receiver3.irq
		.sender_irq    (cpu_d_irq_irq)                   //    sender.irq
	);

endmodule
