library ieee;
use ieee.std_logic_1164.all;

entity ifft_data_gen is
  generic(N: integer range 0 to 511:=80);
  port(rst_n: in std_logic;
       clk: in std_logic;
       din: in std_logic_vector(415 downto 0);
       frame_flag:in std_logic;
       source_data_valid:in std_logic;
       sink_data_valid:out std_logic;
       sop:out std_logic;
       eop:out std_logic;
       dout_real:out std_logic_vector(11 downto 0);
       dout_imag:out std_logic_vector(11 downto 0));
end entity ifft_data_gen ;

architecture rtl of ifft_data_gen is
 signal cnt,cnt1: integer range 0 to 1023;
 type  phase_t is array ( 0 to 415) of std_logic_vector(3 downto 0);
 constant m_phase:phase_t:= (
"0100","1110","1101","1100","0000","0001","0001","1110","1011",
"0100","1110","1010","1000","0011","0011","0000","0110","1111",
"0011","1011","0110","1010","1111","0111","0100","1100","1101",
"1100","0100","0110","1000","0001","0010","1010","1110","0011",
"0000","1110","0010","1100","1000","0101","1000","0000","0110",
"0001","0101","0111","0011","1001","1100","0010","1011","1001",
"0110","0000","1101","0101","1010","1001","1011","1001","0101",
"0011","1010","1011","0010","1111","1100","1100","0111","0011",
"1011","0011","0010","1100","1001","1010","1011","0010","1010",
"0000","0001","0111","0110","0010","0000","0010","0100","0010",
"1001","0010","0011","1000","1101","1011","1111","0101","1000",
"1000","1000","1011","0001","0011","1011","1110","0101","0101",
"1110","0110","1100","1100","1110","0110","1100","1000","0100",
"0000","1100","0111","0000","0000","0011","0111","1011","1111",
"0000","0101","0001","0110","0010","0000","1111","0011","0101",
"1100","1101","0010","0111","0001","0110","1111","0110","1011",
"0101","0001","0001","1111","0000","1000","0001","0100","1111",
"1111","1101","0010","0000","0100","0001","0100","0110","0010",
"1111","0111","1101","0000","0000","0000","0100","0010","1011",
"1011","1010","1110","1001","0000","0001","1111","1011","1001",
"1111","0100","1011","1001","0101","1000","1011","1001","1010",
"0010","0000","1011","0101","1101","0011","0000","1110","0011",
"0001","0110","1100","0100","1000","1111","1010","0010","0010",
"1010","1111","1011","1110","1011","1111","0000","1011","1000",
"1011","1011","0101","0110","1111","0111","0011","0001","1001",
"0001","0101","1100","1000","0011","0101","1011","0000","1101",
"1001","0011","1100","1011","1011","1111","0000","1101","0100",
"1111","0000","0011","1101","0000","1101","0101","1000","1110",
"0100","0011","0000","1010","0110","0001","1011","1010","1010",
"1110","1111","1001","0111","1010","1011","0001","0011","1111",
"0011","1101","1101","1111","1010","0100","1111","0010","1111",
"1111","1011","1011","0000","1010","1010","0000","1111","0000",
"1000","1110","0000","1100","0001","0110","1001","1111","1010",
"0101","1100","0110","0100","0010","1011","1011","1100","0001",
"1001","1100","1111","1010","0011","0101","0000","1001","1010",
"0100","0100","1100","1101","1110","0101","0000","0101","0001",
"1001","1011","0010","1011","0011","1000","0101","1000","1101",
"0001","0011","0101","1110","0101","1000","0011","0100","0001",
"1111","1101","1101","1010","0101","0100","0001","1001","1001",
"1011","0111","0111","0110","0011","0110","0110","1010","1111",
"0100","1000","0100","1011","0111","1100","1110","1010","1100",
"1010","1010","1100","0100","0110","0001","1000","0010","1101",
"1000","1011","1111","0111","0111","0010","0011","0100","0000",
"0000","0010","0111","1011","0111","0010","1011","1101","0001",
"0111","0111","0110","0000","1110","1000","0111","0101","1001",
"1010","0011","1011","0000","0000","1110","1101","1110","1111",
"0001","1001");

 
  
  
  signal pre_phase_s:phase_t;
 signal phase_sub_carrier_s:std_logic_vector(3 downto 0);

 begin

  process(rst_n,clk) is
    
    begin
      if rst_n='0' then
         cnt<=0; 
         sop<='0'; 
         eop<='0';        
      elsif clk'event and clk='1' then
        sink_data_valid<=source_data_valid;
          if source_data_valid='1' then
           if cnt=1023 then
               cnt<=0;
           else
              cnt<=cnt+1;
           end if;
		 case cnt is
           when 1023 =>
            sop<='0'; 
            eop<='1';
           when 0 =>
            sop<='1'; 
            eop<='0';
           when others =>
            sop<='0'; 
            eop<='0';
         end case;
		else 
		     cnt<=0;
		     sop<='0'; 
         eop<='0'; 
			 
		 end if;
      end if;
	  
  end process;


	
 process(rst_n,clk) is
   variable phase_sub_carrier:std_logic_vector(3 downto 0);
   variable pre_phase:phase_t;
    begin
    if rst_n<='0' then
       dout_real<=(others=>'0');
       dout_imag<=(others=>'0');
	     pre_phase:=m_phase;
     elsif clk'event and clk='1' then
       if frame_flag='1' then
		     case cnt is	
		       when N to N+415 => 
		          if din(495-cnt)='0' then
                 pre_phase(cnt-80):=pre_phase(cnt-80);
              else  
                 pre_phase(cnt-80):=not(pre_phase(cnt-80)(3))&pre_phase(cnt-80)(2 downto 0);
			        end if; 

           phase_sub_carrier:=	pre_phase(cnt-80);  
                  
        case phase_sub_carrier is		
					when "0000"=> 
						dout_real<="001111111111";
						dout_imag<="000000000000";
					when "0001"=> 
						dout_real<="001110110001";
						dout_imag<="000110000111";
					when "0010"=> 
						dout_real<="001011010011";
						dout_imag<="001011010011";
					when "0011"=> 
						dout_real<="000110000111";
						dout_imag<="001110110001";
					when "0100"=> 
						dout_real<="000000000000";
						dout_imag<="001111111111";
					when "0101"=> 
						dout_real<="111001111001";
						dout_imag<="001110110001";
					when "0110"=> 
						dout_real<="110100101101";
						dout_imag<="001011010011";
					when "0111"=> 
						dout_real<="110001001111";
						dout_imag<="000110000111";
					when "1000"=> 
						dout_real<="110000000001";
						dout_imag<="000000000000";	
					when "1001"=> 
						dout_real<="110001001111";
						dout_imag<="111001111001";
					when "1010"=> 
						dout_real<="110100101101";
						dout_imag<="110100101101";
					when "1011"=> 
						dout_real<="111001111001";
						dout_imag<="110001001111";
					when "1100"=> 
						dout_real<="000000000000";
						dout_imag<="110000000001";
					when "1101"=> 
						dout_real<="000110000111";
						dout_imag<="110001001111";
					when "1110"=> 
						dout_real<="001011010011";
						dout_imag<="110100101101";
					when "1111"=> 
						dout_real<="001110110001";
						dout_imag<="111001111001";
				   when others => 
						dout_real<=(others=>'0');
						dout_imag<=(others=>'0');
				end case;				
    when others =>
        dout_real<=(others=>'0');
				dout_imag<=(others=>'0');
    end case;
  else
      dout_real<=(others=>'0');
			dout_imag<=(others=>'0');
      pre_phase:=m_phase;
  end if;
 end if;
 pre_phase_s<=pre_phase;
 phase_sub_carrier_s<=phase_sub_carrier;
 end process;


   
  end architecture rtl;
